../005-success-hybrid-abstract/spm.lef