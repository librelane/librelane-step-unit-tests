module xtea (all_done,
    clock,
    mode,
    reset,
    data_in1,
    data_in2,
    data_out1,
    data_out2,
    key_in);
 output all_done;
 input clock;
 input mode;
 input reset;
 input [31:0] data_in1;
 input [31:0] data_in2;
 output [31:0] data_out1;
 output [31:0] data_out2;
 input [127:0] key_in;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire \delta[0] ;
 wire modereg;
 wire \selectslice[0] ;
 wire \selectslice[1] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \state[4] ;
 wire \sum[0] ;
 wire \sum[10] ;
 wire \sum[11] ;
 wire \sum[12] ;
 wire \sum[13] ;
 wire \sum[14] ;
 wire \sum[15] ;
 wire \sum[16] ;
 wire \sum[17] ;
 wire \sum[18] ;
 wire \sum[19] ;
 wire \sum[1] ;
 wire \sum[20] ;
 wire \sum[21] ;
 wire \sum[22] ;
 wire \sum[23] ;
 wire \sum[24] ;
 wire \sum[25] ;
 wire \sum[26] ;
 wire \sum[27] ;
 wire \sum[28] ;
 wire \sum[29] ;
 wire \sum[2] ;
 wire \sum[30] ;
 wire \sum[31] ;
 wire \sum[3] ;
 wire \sum[4] ;
 wire \sum[5] ;
 wire \sum[6] ;
 wire \sum[7] ;
 wire \sum[8] ;
 wire \sum[9] ;
 wire while_flag;
 wire \workunit1[0] ;
 wire \workunit1[10] ;
 wire \workunit1[11] ;
 wire \workunit1[12] ;
 wire \workunit1[13] ;
 wire \workunit1[14] ;
 wire \workunit1[15] ;
 wire \workunit1[16] ;
 wire \workunit1[17] ;
 wire \workunit1[18] ;
 wire \workunit1[19] ;
 wire \workunit1[1] ;
 wire \workunit1[20] ;
 wire \workunit1[21] ;
 wire \workunit1[22] ;
 wire \workunit1[23] ;
 wire \workunit1[24] ;
 wire \workunit1[25] ;
 wire \workunit1[26] ;
 wire \workunit1[27] ;
 wire \workunit1[28] ;
 wire \workunit1[29] ;
 wire \workunit1[2] ;
 wire \workunit1[30] ;
 wire \workunit1[31] ;
 wire \workunit1[3] ;
 wire \workunit1[4] ;
 wire \workunit1[5] ;
 wire \workunit1[6] ;
 wire \workunit1[7] ;
 wire \workunit1[8] ;
 wire \workunit1[9] ;
 wire \workunit2[0] ;
 wire \workunit2[10] ;
 wire \workunit2[11] ;
 wire \workunit2[12] ;
 wire \workunit2[13] ;
 wire \workunit2[14] ;
 wire \workunit2[15] ;
 wire \workunit2[16] ;
 wire \workunit2[17] ;
 wire \workunit2[18] ;
 wire \workunit2[19] ;
 wire \workunit2[1] ;
 wire \workunit2[20] ;
 wire \workunit2[21] ;
 wire \workunit2[22] ;
 wire \workunit2[23] ;
 wire \workunit2[24] ;
 wire \workunit2[25] ;
 wire \workunit2[26] ;
 wire \workunit2[27] ;
 wire \workunit2[28] ;
 wire \workunit2[29] ;
 wire \workunit2[2] ;
 wire \workunit2[30] ;
 wire \workunit2[31] ;
 wire \workunit2[3] ;
 wire \workunit2[4] ;
 wire \workunit2[5] ;
 wire \workunit2[6] ;
 wire \workunit2[7] ;
 wire \workunit2[8] ;
 wire \workunit2[9] ;
 wire \x[0] ;
 wire \x[1] ;
 wire \x[2] ;
 wire \x[3] ;
 wire \x[4] ;
 wire \x[5] ;
 wire \x[6] ;
 wire \x[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire clknet_0_clock;
 wire clknet_4_0_0_clock;
 wire clknet_4_1_0_clock;
 wire clknet_4_2_0_clock;
 wire clknet_4_3_0_clock;
 wire clknet_4_4_0_clock;
 wire clknet_4_5_0_clock;
 wire clknet_4_6_0_clock;
 wire clknet_4_7_0_clock;
 wire clknet_4_8_0_clock;
 wire clknet_4_9_0_clock;
 wire clknet_4_10_0_clock;
 wire clknet_4_11_0_clock;
 wire clknet_4_12_0_clock;
 wire clknet_4_13_0_clock;
 wire clknet_4_14_0_clock;
 wire clknet_4_15_0_clock;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;

 sky130_fd_sc_hd__a211oi_1 _2195_ (.A1(_1666_),
    .A2(_1665_),
    .B1(_1664_),
    .C1(_1619_),
    .Y(_1755_));
 sky130_fd_sc_hd__o21a_1 _2196_ (.A1(_1667_),
    .A2(_1755_),
    .B1(_1717_),
    .X(_1756_));
 sky130_fd_sc_hd__o21ba_1 _2197_ (.A1(\sum[16] ),
    .A2(_1722_),
    .B1_N(_1756_),
    .X(_0273_));
 sky130_fd_sc_hd__nand2_1 _2198_ (.A(\sum[15] ),
    .B(_1725_),
    .Y(_1757_));
 sky130_fd_sc_hd__o21ai_1 _2199_ (.A1(_1656_),
    .A2(_1658_),
    .B1(_1663_),
    .Y(_1758_));
 sky130_fd_sc_hd__nor2_1 _2200_ (.A(_1661_),
    .B(_1758_),
    .Y(_1759_));
 sky130_fd_sc_hd__a211o_1 _2201_ (.A1(_1757_),
    .A2(_1659_),
    .B1(_1759_),
    .C1(_1618_),
    .X(_1760_));
 sky130_fd_sc_hd__o211ai_1 _2202_ (.A1(_1618_),
    .A2(_1759_),
    .B1(_1659_),
    .C1(_1757_),
    .Y(_1761_));
 sky130_fd_sc_hd__a32o_1 _2203_ (.A1(_1729_),
    .A2(_1760_),
    .A3(_1761_),
    .B1(_1742_),
    .B2(\sum[15] ),
    .X(_0272_));
 sky130_fd_sc_hd__nand2_1 _2204_ (.A(_1661_),
    .B(_1758_),
    .Y(_1762_));
 sky130_fd_sc_hd__nor2_1 _2205_ (.A(_1708_),
    .B(_1759_),
    .Y(_1763_));
 sky130_fd_sc_hd__a22o_1 _2206_ (.A1(\sum[14] ),
    .A2(_1742_),
    .B1(_1762_),
    .B2(_1763_),
    .X(_0271_));
 sky130_fd_sc_hd__a21o_1 _2207_ (.A1(net379),
    .A2(_1704_),
    .B1(_1656_),
    .X(_1764_));
 sky130_fd_sc_hd__a21boi_1 _2208_ (.A1(_1663_),
    .A2(_1657_),
    .B1_N(_1764_),
    .Y(_1765_));
 sky130_fd_sc_hd__and3b_1 _2209_ (.A_N(_1764_),
    .B(_1657_),
    .C(_1663_),
    .X(_1766_));
 sky130_fd_sc_hd__o32a_1 _2210_ (.A1(_1708_),
    .A2(_1765_),
    .A3(_1766_),
    .B1(_1739_),
    .B2(net592),
    .X(_0270_));
 sky130_fd_sc_hd__or2_1 _2211_ (.A(_1621_),
    .B(_1650_),
    .X(_1767_));
 sky130_fd_sc_hd__a211o_1 _2212_ (.A1(_1655_),
    .A2(_1767_),
    .B1(_1654_),
    .C1(_1620_),
    .X(_1768_));
 sky130_fd_sc_hd__and2b_1 _2213_ (.A_N(_1656_),
    .B(_1768_),
    .X(_1769_));
 sky130_fd_sc_hd__o22a_1 _2214_ (.A1(net379),
    .A2(_1598_),
    .B1(_1769_),
    .B2(_1711_),
    .X(_0269_));
 sky130_fd_sc_hd__nand2_1 _2215_ (.A(net380),
    .B(_1704_),
    .Y(_1770_));
 sky130_fd_sc_hd__nand2_1 _2216_ (.A(_1655_),
    .B(_1770_),
    .Y(_1771_));
 sky130_fd_sc_hd__xnor2_1 _2217_ (.A(_1767_),
    .B(_1771_),
    .Y(_1772_));
 sky130_fd_sc_hd__a22o_1 _2218_ (.A1(net381),
    .A2(_1742_),
    .B1(_1772_),
    .B2(_1729_),
    .X(_0268_));
 sky130_fd_sc_hd__nand2_1 _2219_ (.A(_1624_),
    .B(_1649_),
    .Y(_1773_));
 sky130_fd_sc_hd__xnor2_1 _2220_ (.A(_1623_),
    .B(_1773_),
    .Y(_1774_));
 sky130_fd_sc_hd__o2bb2a_1 _2221_ (.A1_N(_1718_),
    .A2_N(_1774_),
    .B1(_1722_),
    .B2(\sum[10] ),
    .X(_0267_));
 sky130_fd_sc_hd__nor2_1 _2222_ (.A(net382),
    .B(_1725_),
    .Y(_1775_));
 sky130_fd_sc_hd__a21o_1 _2223_ (.A1(_1645_),
    .A2(_1646_),
    .B1(_1648_),
    .X(_1776_));
 sky130_fd_sc_hd__nor3_1 _2224_ (.A(_1775_),
    .B(_1647_),
    .C(_1776_),
    .Y(_1777_));
 sky130_fd_sc_hd__o21a_1 _2225_ (.A1(_1775_),
    .A2(_1647_),
    .B1(_1776_),
    .X(_1778_));
 sky130_fd_sc_hd__o32a_1 _2226_ (.A1(_1708_),
    .A2(_1777_),
    .A3(_1778_),
    .B1(_1739_),
    .B2(net382),
    .X(_0266_));
 sky130_fd_sc_hd__or2b_1 _2227_ (.A(_1648_),
    .B_N(_1646_),
    .X(_1779_));
 sky130_fd_sc_hd__xnor2_1 _2228_ (.A(_1645_),
    .B(_1779_),
    .Y(_1780_));
 sky130_fd_sc_hd__o22a_1 _2229_ (.A1(net594),
    .A2(_1598_),
    .B1(_1780_),
    .B2(_1711_),
    .X(_0265_));
 sky130_fd_sc_hd__nand3_1 _2230_ (.A(_1644_),
    .B(_1625_),
    .C(_1643_),
    .Y(_1781_));
 sky130_fd_sc_hd__a21o_1 _2231_ (.A1(_1644_),
    .A2(_1625_),
    .B1(_1643_),
    .X(_1782_));
 sky130_fd_sc_hd__a32o_1 _2232_ (.A1(_1729_),
    .A2(_1781_),
    .A3(_1782_),
    .B1(_1742_),
    .B2(\sum[7] ),
    .X(_0264_));
 sky130_fd_sc_hd__and2_1 _2233_ (.A(net383),
    .B(_1725_),
    .X(_1783_));
 sky130_fd_sc_hd__nor4_1 _2234_ (.A(_1783_),
    .B(_1626_),
    .C(_1627_),
    .D(_1641_),
    .Y(_1784_));
 sky130_fd_sc_hd__o22a_1 _2235_ (.A1(_1783_),
    .A2(_1626_),
    .B1(_1627_),
    .B2(_1641_),
    .X(_1785_));
 sky130_fd_sc_hd__nor2_1 _2236_ (.A(_1784_),
    .B(_1785_),
    .Y(_1786_));
 sky130_fd_sc_hd__a22o_1 _2237_ (.A1(net383),
    .A2(_1714_),
    .B1(_1786_),
    .B2(_1718_),
    .X(_0263_));
 sky130_fd_sc_hd__and2b_1 _2238_ (.A_N(_1627_),
    .B(_1641_),
    .X(_1787_));
 sky130_fd_sc_hd__and2_1 _2239_ (.A(_1636_),
    .B(_1639_),
    .X(_1788_));
 sky130_fd_sc_hd__o22a_1 _2240_ (.A1(_1627_),
    .A2(_1640_),
    .B1(_1637_),
    .B2(_1788_),
    .X(_1789_));
 sky130_fd_sc_hd__o32a_1 _2241_ (.A1(_1708_),
    .A2(_1787_),
    .A3(_1789_),
    .B1(_1739_),
    .B2(\sum[5] ),
    .X(_0262_));
 sky130_fd_sc_hd__or2_1 _2242_ (.A(_1636_),
    .B(_1639_),
    .X(_1790_));
 sky130_fd_sc_hd__nor2_1 _2243_ (.A(_1707_),
    .B(_1788_),
    .Y(_1791_));
 sky130_fd_sc_hd__a22o_1 _2244_ (.A1(\sum[4] ),
    .A2(_1714_),
    .B1(_1790_),
    .B2(_1791_),
    .X(_0261_));
 sky130_fd_sc_hd__and3_1 _2245_ (.A(_1635_),
    .B(_1628_),
    .C(_1634_),
    .X(_1792_));
 sky130_fd_sc_hd__inv_2 _2246_ (.A(_1792_),
    .Y(_1793_));
 sky130_fd_sc_hd__a21o_1 _2247_ (.A1(_1635_),
    .A2(_1628_),
    .B1(_1634_),
    .X(_1794_));
 sky130_fd_sc_hd__a32o_1 _2248_ (.A1(_1729_),
    .A2(_1793_),
    .A3(_1794_),
    .B1(_1742_),
    .B2(net593),
    .X(_0260_));
 sky130_fd_sc_hd__or2b_1 _2249_ (.A(_1633_),
    .B_N(_1632_),
    .X(_1795_));
 sky130_fd_sc_hd__xnor2_1 _2250_ (.A(_1631_),
    .B(_1795_),
    .Y(_1796_));
 sky130_fd_sc_hd__a22o_1 _2251_ (.A1(\sum[2] ),
    .A2(_1714_),
    .B1(_1796_),
    .B2(_1718_),
    .X(_0259_));
 sky130_fd_sc_hd__nand2_1 _2252_ (.A(net384),
    .B(_1725_),
    .Y(_1797_));
 sky130_fd_sc_hd__and4_1 _2253_ (.A(net385),
    .B(net398),
    .C(_1797_),
    .D(_1629_),
    .X(_1798_));
 sky130_fd_sc_hd__inv_2 _2254_ (.A(_1798_),
    .Y(_1799_));
 sky130_fd_sc_hd__a22o_1 _2255_ (.A1(net385),
    .A2(net398),
    .B1(_1797_),
    .B2(_1629_),
    .X(_1800_));
 sky130_fd_sc_hd__a32o_1 _2256_ (.A1(_1729_),
    .A2(_1799_),
    .A3(_1800_),
    .B1(_1713_),
    .B2(net591),
    .X(_0258_));
 sky130_fd_sc_hd__a21o_1 _2257_ (.A1(net385),
    .A2(net398),
    .B1(_1707_),
    .X(_1801_));
 sky130_fd_sc_hd__a21oi_1 _2258_ (.A1(net399),
    .A2(_1597_),
    .B1(net385),
    .Y(_1802_));
 sky130_fd_sc_hd__a21oi_1 _2259_ (.A1(_1739_),
    .A2(_1801_),
    .B1(_1802_),
    .Y(_0257_));
 sky130_fd_sc_hd__nor2_1 _2260_ (.A(net265),
    .B(_0999_),
    .Y(_1803_));
 sky130_fd_sc_hd__o211a_1 _2261_ (.A1(_0669_),
    .A2(_1803_),
    .B1(\x[1] ),
    .C1(\x[0] ),
    .X(_1804_));
 sky130_fd_sc_hd__and2_1 _2262_ (.A(\x[2] ),
    .B(_1804_),
    .X(_1805_));
 sky130_fd_sc_hd__and3_1 _2263_ (.A(\x[4] ),
    .B(\x[3] ),
    .C(_1805_),
    .X(_1806_));
 sky130_fd_sc_hd__and2_1 _2264_ (.A(\x[5] ),
    .B(_1806_),
    .X(_1807_));
 sky130_fd_sc_hd__nand2_1 _2265_ (.A(\x[6] ),
    .B(_1807_),
    .Y(_1808_));
 sky130_fd_sc_hd__xnor2_1 _2266_ (.A(net585),
    .B(_1808_),
    .Y(_0256_));
 sky130_fd_sc_hd__or2_1 _2267_ (.A(\x[6] ),
    .B(_1807_),
    .X(_1809_));
 sky130_fd_sc_hd__and2_1 _2268_ (.A(_1808_),
    .B(_1809_),
    .X(_1810_));
 sky130_fd_sc_hd__clkbuf_1 _2269_ (.A(_1810_),
    .X(_0255_));
 sky130_fd_sc_hd__nor2_1 _2270_ (.A(net590),
    .B(_1806_),
    .Y(_1811_));
 sky130_fd_sc_hd__nor2_1 _2271_ (.A(_1807_),
    .B(_1811_),
    .Y(_0254_));
 sky130_fd_sc_hd__a21oi_1 _2272_ (.A1(net587),
    .A2(_1805_),
    .B1(net589),
    .Y(_1812_));
 sky130_fd_sc_hd__nor2_1 _2273_ (.A(_1806_),
    .B(_1812_),
    .Y(_0253_));
 sky130_fd_sc_hd__xor2_1 _2274_ (.A(net587),
    .B(_1805_),
    .X(_0252_));
 sky130_fd_sc_hd__nor2_1 _2275_ (.A(net588),
    .B(_1804_),
    .Y(_1813_));
 sky130_fd_sc_hd__nor2_1 _2276_ (.A(_1805_),
    .B(_1813_),
    .Y(_0251_));
 sky130_fd_sc_hd__o21ai_1 _2277_ (.A1(_0669_),
    .A2(_1803_),
    .B1(\x[0] ),
    .Y(_1814_));
 sky130_fd_sc_hd__xnor2_1 _2278_ (.A(net586),
    .B(_1814_),
    .Y(_0250_));
 sky130_fd_sc_hd__or3_1 _2279_ (.A(\x[0] ),
    .B(_0669_),
    .C(_1803_),
    .X(_1815_));
 sky130_fd_sc_hd__and2_1 _2280_ (.A(_1814_),
    .B(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__clkbuf_1 _2281_ (.A(_1816_),
    .X(_0249_));
 sky130_fd_sc_hd__or3_2 _2282_ (.A(\state[4] ),
    .B(\state[0] ),
    .C(_0998_),
    .X(_1817_));
 sky130_fd_sc_hd__nand2_1 _2283_ (.A(net263),
    .B(_0871_),
    .Y(_1818_));
 sky130_fd_sc_hd__inv_2 _2284_ (.A(_1817_),
    .Y(_1819_));
 sky130_fd_sc_hd__a32o_1 _2285_ (.A1(net379),
    .A2(net263),
    .A3(_0871_),
    .B1(_1819_),
    .B2(\sum[1] ),
    .X(_1820_));
 sky130_fd_sc_hd__a31o_1 _2286_ (.A1(net389),
    .A2(_1817_),
    .A3(_1818_),
    .B1(_1820_),
    .X(_0248_));
 sky130_fd_sc_hd__nand2_1 _2287_ (.A(_1817_),
    .B(_1818_),
    .Y(_1821_));
 sky130_fd_sc_hd__or2_1 _2288_ (.A(net395),
    .B(_1821_),
    .X(_1822_));
 sky130_fd_sc_hd__o221a_1 _2289_ (.A1(\sum[0] ),
    .A2(_1817_),
    .B1(_1818_),
    .B2(net381),
    .C1(_1822_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _2290_ (.A0(modereg),
    .A1(net533),
    .S(_0893_),
    .X(_1823_));
 sky130_fd_sc_hd__clkbuf_1 _2291_ (.A(_1823_),
    .X(_0246_));
 sky130_fd_sc_hd__nor3_1 _2292_ (.A(\x[7] ),
    .B(\x[6] ),
    .C(\x[5] ),
    .Y(_1824_));
 sky130_fd_sc_hd__and3_1 _2293_ (.A(_0867_),
    .B(_0769_),
    .C(_0512_),
    .X(_1825_));
 sky130_fd_sc_hd__mux2_1 _2294_ (.A0(while_flag),
    .A1(_1824_),
    .S(_1825_),
    .X(_1826_));
 sky130_fd_sc_hd__clkbuf_1 _2295_ (.A(_1826_),
    .X(_0245_));
 sky130_fd_sc_hd__and4_1 _2296_ (.A(\state[4] ),
    .B(_0997_),
    .C(_0867_),
    .D(_0769_),
    .X(_1827_));
 sky130_fd_sc_hd__and2_1 _2297_ (.A(\state[0] ),
    .B(_1827_),
    .X(_1828_));
 sky130_fd_sc_hd__or2_1 _2298_ (.A(net195),
    .B(_1828_),
    .X(_1829_));
 sky130_fd_sc_hd__clkbuf_1 _2299_ (.A(_1829_),
    .X(_0244_));
 sky130_fd_sc_hd__or3b_1 _2300_ (.A(_0867_),
    .B(net261),
    .C_N(_1922_),
    .X(_1830_));
 sky130_fd_sc_hd__nor2_1 _2301_ (.A(net264),
    .B(_1830_),
    .Y(_1831_));
 sky130_fd_sc_hd__and3_1 _2302_ (.A(net262),
    .B(net261),
    .C(_1594_),
    .X(_1832_));
 sky130_fd_sc_hd__a211o_1 _2303_ (.A1(_0512_),
    .A2(_0998_),
    .B1(_1831_),
    .C1(_1832_),
    .X(_1833_));
 sky130_fd_sc_hd__nor3_1 _2304_ (.A(_1821_),
    .B(_1828_),
    .C(_1833_),
    .Y(_1834_));
 sky130_fd_sc_hd__o211a_2 _2305_ (.A1(net262),
    .A2(_0870_),
    .B1(_1596_),
    .C1(_1834_),
    .X(_1835_));
 sky130_fd_sc_hd__clkbuf_4 _2306_ (.A(_1835_),
    .X(_1836_));
 sky130_fd_sc_hd__clkbuf_4 _2307_ (.A(_1836_),
    .X(_1837_));
 sky130_fd_sc_hd__mux2_1 _2308_ (.A0(net252),
    .A1(\workunit2[31] ),
    .S(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__clkbuf_1 _2309_ (.A(_1838_),
    .X(_0243_));
 sky130_fd_sc_hd__clkbuf_4 _2310_ (.A(_1835_),
    .X(_1839_));
 sky130_fd_sc_hd__buf_2 _2311_ (.A(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__mux2_1 _2312_ (.A0(net251),
    .A1(net266),
    .S(_1840_),
    .X(_1841_));
 sky130_fd_sc_hd__clkbuf_1 _2313_ (.A(_1841_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _2314_ (.A0(net249),
    .A1(\workunit2[29] ),
    .S(_1840_),
    .X(_1842_));
 sky130_fd_sc_hd__clkbuf_1 _2315_ (.A(_1842_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _2316_ (.A0(net248),
    .A1(\workunit2[28] ),
    .S(_1840_),
    .X(_1843_));
 sky130_fd_sc_hd__clkbuf_1 _2317_ (.A(_1843_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _2318_ (.A0(net247),
    .A1(net270),
    .S(_1840_),
    .X(_1844_));
 sky130_fd_sc_hd__clkbuf_1 _2319_ (.A(_1844_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _2320_ (.A0(net246),
    .A1(net272),
    .S(_1840_),
    .X(_1845_));
 sky130_fd_sc_hd__clkbuf_1 _2321_ (.A(_1845_),
    .X(_0238_));
 sky130_fd_sc_hd__clkbuf_2 _2322_ (.A(_1839_),
    .X(_1846_));
 sky130_fd_sc_hd__mux2_1 _2323_ (.A0(net245),
    .A1(net274),
    .S(_1846_),
    .X(_1847_));
 sky130_fd_sc_hd__clkbuf_1 _2324_ (.A(_1847_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _2325_ (.A0(net244),
    .A1(net277),
    .S(_1846_),
    .X(_1848_));
 sky130_fd_sc_hd__clkbuf_1 _2326_ (.A(_1848_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _2327_ (.A0(net243),
    .A1(net279),
    .S(_1846_),
    .X(_1849_));
 sky130_fd_sc_hd__clkbuf_1 _2328_ (.A(_1849_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _2329_ (.A0(net242),
    .A1(net281),
    .S(_1846_),
    .X(_1850_));
 sky130_fd_sc_hd__clkbuf_1 _2330_ (.A(_1850_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _2331_ (.A0(net241),
    .A1(net282),
    .S(_1846_),
    .X(_1851_));
 sky130_fd_sc_hd__clkbuf_1 _2332_ (.A(_1851_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _2333_ (.A0(net240),
    .A1(net285),
    .S(_1846_),
    .X(_1852_));
 sky130_fd_sc_hd__clkbuf_1 _2334_ (.A(_1852_),
    .X(_0232_));
 sky130_fd_sc_hd__clkbuf_2 _2335_ (.A(_1836_),
    .X(_1853_));
 sky130_fd_sc_hd__mux2_1 _2336_ (.A0(net238),
    .A1(net288),
    .S(_1853_),
    .X(_1854_));
 sky130_fd_sc_hd__clkbuf_1 _2337_ (.A(_1854_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _2338_ (.A0(net237),
    .A1(net290),
    .S(_1853_),
    .X(_1855_));
 sky130_fd_sc_hd__clkbuf_1 _2339_ (.A(_1855_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _2340_ (.A0(net236),
    .A1(net292),
    .S(_1853_),
    .X(_1856_));
 sky130_fd_sc_hd__clkbuf_1 _2341_ (.A(_1856_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _2342_ (.A0(net235),
    .A1(net294),
    .S(_1853_),
    .X(_1857_));
 sky130_fd_sc_hd__clkbuf_1 _2343_ (.A(_1857_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _2344_ (.A0(net234),
    .A1(\workunit2[15] ),
    .S(_1853_),
    .X(_1858_));
 sky130_fd_sc_hd__clkbuf_1 _2345_ (.A(_1858_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _2346_ (.A0(net233),
    .A1(net298),
    .S(_1853_),
    .X(_1859_));
 sky130_fd_sc_hd__clkbuf_1 _2347_ (.A(_1859_),
    .X(_0226_));
 sky130_fd_sc_hd__clkbuf_2 _2348_ (.A(_1836_),
    .X(_1860_));
 sky130_fd_sc_hd__mux2_1 _2349_ (.A0(net232),
    .A1(net300),
    .S(_1860_),
    .X(_1861_));
 sky130_fd_sc_hd__clkbuf_1 _2350_ (.A(_1861_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _2351_ (.A0(net231),
    .A1(net302),
    .S(_1860_),
    .X(_1862_));
 sky130_fd_sc_hd__clkbuf_1 _2352_ (.A(_1862_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _2353_ (.A0(net230),
    .A1(net304),
    .S(_1860_),
    .X(_1863_));
 sky130_fd_sc_hd__clkbuf_1 _2354_ (.A(_1863_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _2355_ (.A0(net229),
    .A1(net306),
    .S(_1860_),
    .X(_1864_));
 sky130_fd_sc_hd__clkbuf_1 _2356_ (.A(_1864_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _2357_ (.A0(net259),
    .A1(net308),
    .S(_1860_),
    .X(_1865_));
 sky130_fd_sc_hd__clkbuf_1 _2358_ (.A(_1865_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _2359_ (.A0(net258),
    .A1(net310),
    .S(_1860_),
    .X(_1866_));
 sky130_fd_sc_hd__clkbuf_1 _2360_ (.A(_1866_),
    .X(_0220_));
 sky130_fd_sc_hd__clkbuf_2 _2361_ (.A(_1836_),
    .X(_1867_));
 sky130_fd_sc_hd__mux2_1 _2362_ (.A0(net257),
    .A1(net311),
    .S(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__clkbuf_1 _2363_ (.A(_1868_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _2364_ (.A0(net256),
    .A1(net313),
    .S(_1867_),
    .X(_1869_));
 sky130_fd_sc_hd__clkbuf_1 _2365_ (.A(_1869_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _2366_ (.A0(net255),
    .A1(net316),
    .S(_1867_),
    .X(_1870_));
 sky130_fd_sc_hd__clkbuf_1 _2367_ (.A(_1870_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _2368_ (.A0(net254),
    .A1(\workunit2[4] ),
    .S(_1867_),
    .X(_1871_));
 sky130_fd_sc_hd__clkbuf_1 _2369_ (.A(_1871_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _2370_ (.A0(net253),
    .A1(\workunit2[3] ),
    .S(_1867_),
    .X(_1872_));
 sky130_fd_sc_hd__clkbuf_1 _2371_ (.A(_1872_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _2372_ (.A0(net250),
    .A1(net320),
    .S(_1867_),
    .X(_1873_));
 sky130_fd_sc_hd__clkbuf_1 _2373_ (.A(_1873_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _2374_ (.A0(net239),
    .A1(net321),
    .S(_1837_),
    .X(_1874_));
 sky130_fd_sc_hd__clkbuf_1 _2375_ (.A(_1874_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _2376_ (.A0(net228),
    .A1(net322),
    .S(_1837_),
    .X(_1875_));
 sky130_fd_sc_hd__clkbuf_1 _2377_ (.A(_1875_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _2378_ (.A0(net220),
    .A1(\workunit1[31] ),
    .S(_1839_),
    .X(_1876_));
 sky130_fd_sc_hd__clkbuf_1 _2379_ (.A(_1876_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _2380_ (.A0(net219),
    .A1(\workunit1[30] ),
    .S(_1837_),
    .X(_1877_));
 sky130_fd_sc_hd__clkbuf_1 _2381_ (.A(_1877_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _2382_ (.A0(net217),
    .A1(\workunit1[29] ),
    .S(_1837_),
    .X(_1878_));
 sky130_fd_sc_hd__clkbuf_1 _2383_ (.A(_1878_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _2384_ (.A0(net216),
    .A1(\workunit1[28] ),
    .S(_1837_),
    .X(_1879_));
 sky130_fd_sc_hd__clkbuf_1 _2385_ (.A(_1879_),
    .X(_0208_));
 sky130_fd_sc_hd__clkbuf_2 _2386_ (.A(_1836_),
    .X(_1880_));
 sky130_fd_sc_hd__mux2_1 _2387_ (.A0(net215),
    .A1(net326),
    .S(_1880_),
    .X(_1881_));
 sky130_fd_sc_hd__clkbuf_1 _2388_ (.A(_1881_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _2389_ (.A0(net214),
    .A1(net329),
    .S(_1880_),
    .X(_1882_));
 sky130_fd_sc_hd__clkbuf_1 _2390_ (.A(_1882_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _2391_ (.A0(net213),
    .A1(net331),
    .S(_1880_),
    .X(_1883_));
 sky130_fd_sc_hd__clkbuf_1 _2392_ (.A(_1883_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _2393_ (.A0(net212),
    .A1(net333),
    .S(_1880_),
    .X(_1884_));
 sky130_fd_sc_hd__clkbuf_1 _2394_ (.A(_1884_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _2395_ (.A0(net211),
    .A1(net334),
    .S(_1880_),
    .X(_1885_));
 sky130_fd_sc_hd__clkbuf_1 _2396_ (.A(_1885_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _2397_ (.A0(net210),
    .A1(net337),
    .S(_1880_),
    .X(_1886_));
 sky130_fd_sc_hd__clkbuf_1 _2398_ (.A(_1886_),
    .X(_0202_));
 sky130_fd_sc_hd__clkbuf_2 _2399_ (.A(_1836_),
    .X(_1887_));
 sky130_fd_sc_hd__mux2_1 _2400_ (.A0(net209),
    .A1(net338),
    .S(_1887_),
    .X(_1888_));
 sky130_fd_sc_hd__clkbuf_1 _2401_ (.A(_1888_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _2402_ (.A0(net208),
    .A1(net340),
    .S(_1887_),
    .X(_1889_));
 sky130_fd_sc_hd__clkbuf_1 _2403_ (.A(_1889_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _2404_ (.A0(net206),
    .A1(net343),
    .S(_1887_),
    .X(_1890_));
 sky130_fd_sc_hd__clkbuf_1 _2405_ (.A(_1890_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _2406_ (.A0(net205),
    .A1(net345),
    .S(_1887_),
    .X(_1891_));
 sky130_fd_sc_hd__clkbuf_1 _2407_ (.A(_1891_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _2408_ (.A0(net204),
    .A1(net347),
    .S(_1887_),
    .X(_1892_));
 sky130_fd_sc_hd__clkbuf_1 _2409_ (.A(_1892_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _2410_ (.A0(net203),
    .A1(net349),
    .S(_1887_),
    .X(_1893_));
 sky130_fd_sc_hd__clkbuf_1 _2411_ (.A(_1893_),
    .X(_0196_));
 sky130_fd_sc_hd__clkbuf_2 _2412_ (.A(_1835_),
    .X(_1894_));
 sky130_fd_sc_hd__mux2_1 _2413_ (.A0(net202),
    .A1(net351),
    .S(_1894_),
    .X(_1895_));
 sky130_fd_sc_hd__clkbuf_1 _2414_ (.A(_1895_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _2415_ (.A0(net201),
    .A1(net353),
    .S(_1894_),
    .X(_1896_));
 sky130_fd_sc_hd__clkbuf_1 _2416_ (.A(_1896_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _2417_ (.A0(net200),
    .A1(net355),
    .S(_1894_),
    .X(_1897_));
 sky130_fd_sc_hd__clkbuf_1 _2418_ (.A(_1897_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _2419_ (.A0(net199),
    .A1(net357),
    .S(_1894_),
    .X(_1898_));
 sky130_fd_sc_hd__clkbuf_1 _2420_ (.A(_1898_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _2421_ (.A0(net198),
    .A1(net358),
    .S(_1894_),
    .X(_1899_));
 sky130_fd_sc_hd__clkbuf_1 _2422_ (.A(_1899_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _2423_ (.A0(net197),
    .A1(net361),
    .S(_1894_),
    .X(_1900_));
 sky130_fd_sc_hd__clkbuf_1 _2424_ (.A(_1900_),
    .X(_0190_));
 sky130_fd_sc_hd__clkbuf_2 _2425_ (.A(_1835_),
    .X(_1901_));
 sky130_fd_sc_hd__mux2_1 _2426_ (.A0(net227),
    .A1(net363),
    .S(_1901_),
    .X(_1902_));
 sky130_fd_sc_hd__clkbuf_1 _2427_ (.A(_1902_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _2428_ (.A0(net226),
    .A1(net364),
    .S(_1901_),
    .X(_1903_));
 sky130_fd_sc_hd__clkbuf_1 _2429_ (.A(_1903_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _2430_ (.A0(net225),
    .A1(net366),
    .S(_1901_),
    .X(_1904_));
 sky130_fd_sc_hd__clkbuf_1 _2431_ (.A(_1904_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _2432_ (.A0(net224),
    .A1(net368),
    .S(_1901_),
    .X(_1905_));
 sky130_fd_sc_hd__clkbuf_1 _2433_ (.A(_1905_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _2434_ (.A0(net223),
    .A1(net371),
    .S(_1901_),
    .X(_1906_));
 sky130_fd_sc_hd__clkbuf_1 _2435_ (.A(_1906_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _2436_ (.A0(net222),
    .A1(net372),
    .S(_1901_),
    .X(_1907_));
 sky130_fd_sc_hd__clkbuf_1 _2437_ (.A(_1907_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _2438_ (.A0(net221),
    .A1(net373),
    .S(_1839_),
    .X(_1908_));
 sky130_fd_sc_hd__clkbuf_1 _2439_ (.A(_1908_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _2440_ (.A0(net218),
    .A1(net374),
    .S(_1839_),
    .X(_1909_));
 sky130_fd_sc_hd__clkbuf_1 _2441_ (.A(_1909_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _2442_ (.A0(net207),
    .A1(net375),
    .S(_1839_),
    .X(_1910_));
 sky130_fd_sc_hd__clkbuf_1 _2443_ (.A(_1910_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _2444_ (.A0(net196),
    .A1(\workunit1[0] ),
    .S(_1840_),
    .X(_1911_));
 sky130_fd_sc_hd__clkbuf_1 _2445_ (.A(_1911_),
    .X(_0180_));
 sky130_fd_sc_hd__nand2_1 _2446_ (.A(_1600_),
    .B(_1542_),
    .Y(_0179_));
 sky130_fd_sc_hd__a21oi_1 _2447_ (.A1(modereg),
    .A2(_0997_),
    .B1(_1830_),
    .Y(_1912_));
 sky130_fd_sc_hd__a2111o_1 _2448_ (.A1(_0867_),
    .A2(_1922_),
    .B1(_1593_),
    .C1(_1827_),
    .D1(_1912_),
    .X(_2190_));
 sky130_fd_sc_hd__or2_1 _2449_ (.A(_0997_),
    .B(_0870_),
    .X(_1913_));
 sky130_fd_sc_hd__or4_1 _2450_ (.A(while_flag),
    .B(net263),
    .C(\state[3] ),
    .D(_1913_),
    .X(_1914_));
 sky130_fd_sc_hd__a21bo_1 _2451_ (.A1(modereg),
    .A2(_1831_),
    .B1_N(_1914_),
    .X(_1915_));
 sky130_fd_sc_hd__or3_1 _2452_ (.A(_0512_),
    .B(_0871_),
    .C(_1915_),
    .X(_1916_));
 sky130_fd_sc_hd__clkbuf_1 _2453_ (.A(_1916_),
    .X(_2191_));
 sky130_fd_sc_hd__o21ai_1 _2454_ (.A1(net263),
    .A2(_1913_),
    .B1(_1818_),
    .Y(_1917_));
 sky130_fd_sc_hd__or3_1 _2455_ (.A(_1593_),
    .B(_1912_),
    .C(_1917_),
    .X(_1918_));
 sky130_fd_sc_hd__clkbuf_1 _2456_ (.A(_1918_),
    .X(_2192_));
 sky130_fd_sc_hd__nand2_1 _2457_ (.A(_1592_),
    .B(_1817_),
    .Y(_1919_));
 sky130_fd_sc_hd__or4_1 _2458_ (.A(_1002_),
    .B(_1595_),
    .C(_1915_),
    .D(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__clkbuf_1 _2459_ (.A(_1920_),
    .X(_2193_));
 sky130_fd_sc_hd__or2_1 _2460_ (.A(_1827_),
    .B(_1832_),
    .X(_1921_));
 sky130_fd_sc_hd__clkbuf_1 _2461_ (.A(_1921_),
    .X(_2194_));
 sky130_fd_sc_hd__inv_2 _2462_ (.A(net406),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _2463_ (.A(net433),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _2464_ (.A(net405),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _2465_ (.A(net405),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _2466_ (.A(net405),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _2467_ (.A(net406),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _2468_ (.A(net400),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _2469_ (.A(net406),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _2470_ (.A(net406),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _2471_ (.A(net406),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _2472_ (.A(net400),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _2473_ (.A(net422),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _2474_ (.A(net422),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _2475_ (.A(net422),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _2476_ (.A(net424),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _2477_ (.A(net425),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _2478_ (.A(net424),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _2479_ (.A(net427),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _2480_ (.A(net428),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _2481_ (.A(net427),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _2482_ (.A(net427),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _2483_ (.A(net428),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _2484_ (.A(net428),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _2485_ (.A(net430),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _2486_ (.A(net430),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _2487_ (.A(net430),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _2488_ (.A(net430),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _2489_ (.A(net430),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _2490_ (.A(net430),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _2491_ (.A(net433),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _2492_ (.A(net433),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _2493_ (.A(net433),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _2494_ (.A(net433),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _2495_ (.A(net419),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _2496_ (.A(net419),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _2497_ (.A(net414),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _2498_ (.A(net415),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _2499_ (.A(net415),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _2500_ (.A(net414),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _2501_ (.A(net415),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _2502_ (.A(net414),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _2503_ (.A(net414),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _2504_ (.A(net415),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _2505_ (.A(net415),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _2506_ (.A(net415),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _2507_ (.A(net416),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _2508_ (.A(net416),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _2509_ (.A(net435),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _2510_ (.A(net435),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _2511_ (.A(net435),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _2512_ (.A(net435),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _2513_ (.A(net437),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _2514_ (.A(net437),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _2515_ (.A(net443),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _2516_ (.A(net440),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _2517_ (.A(net440),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _2518_ (.A(net440),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _2519_ (.A(net441),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _2520_ (.A(net441),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _2521_ (.A(net442),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _2522_ (.A(net444),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _2523_ (.A(net442),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _2524_ (.A(net441),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _2525_ (.A(net444),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _2526_ (.A(net444),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _2527_ (.A(net400),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _2528_ (.A(net407),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _2529_ (.A(net400),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _2530_ (.A(net402),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _2531_ (.A(net402),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _2532_ (.A(net407),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _2533_ (.A(net407),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _2534_ (.A(net408),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _2535_ (.A(net408),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _2536_ (.A(net419),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _2537_ (.A(net419),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _2538_ (.A(net419),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _2539_ (.A(net419),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _2540_ (.A(net402),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _2541_ (.A(net402),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _2542_ (.A(net400),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _2543_ (.A(net402),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _2544_ (.A(net401),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _2545_ (.A(net401),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _2546_ (.A(net401),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _2547_ (.A(net403),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _2548_ (.A(net403),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _2549_ (.A(net403),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _2550_ (.A(net403),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _2551_ (.A(net402),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _2552_ (.A(net404),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _2553_ (.A(net410),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _2554_ (.A(net403),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _2555_ (.A(net410),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _2556_ (.A(net410),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _2557_ (.A(net410),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _2558_ (.A(net410),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _2559_ (.A(net410),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _2560_ (.A(net413),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _2561_ (.A(net413),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _2562_ (.A(net411),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _2563_ (.A(net411),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _2564_ (.A(net411),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _2565_ (.A(net411),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _2566_ (.A(net412),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _2567_ (.A(net412),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _2568_ (.A(net412),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _2569_ (.A(net412),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _2570_ (.A(net411),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _2571_ (.A(net411),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _2572_ (.A(net406),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _2573_ (.A(net409),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _2574_ (.A(net405),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _2575_ (.A(net405),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _2576_ (.A(net405),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _2577_ (.A(net400),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _2578_ (.A(net422),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _2579_ (.A(net422),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _2580_ (.A(net422),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _2581_ (.A(net426),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _2582_ (.A(net423),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _2583_ (.A(net423),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _2584_ (.A(net424),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _2585_ (.A(net424),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _2586_ (.A(net425),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _2587_ (.A(net424),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _2588_ (.A(net425),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _2589_ (.A(net424),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _2590_ (.A(net425),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _2591_ (.A(net429),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _2592_ (.A(net427),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _2593_ (.A(net425),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _2594_ (.A(net428),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _2595_ (.A(net427),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _2596_ (.A(net429),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _2597_ (.A(net431),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _2598_ (.A(net427),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _2599_ (.A(net431),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _2600_ (.A(net429),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _2601_ (.A(net431),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _2602_ (.A(net434),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _2603_ (.A(net431),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _2604_ (.A(net414),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _2605_ (.A(net418),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _2606_ (.A(net414),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _2607_ (.A(net417),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _2608_ (.A(net417),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _2609_ (.A(net435),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _2610_ (.A(net416),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _2611_ (.A(net436),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _2612_ (.A(net436),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _2613_ (.A(net435),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _2614_ (.A(net436),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _2615_ (.A(net439),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _2616_ (.A(net436),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _2617_ (.A(net436),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _2618_ (.A(net437),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _2619_ (.A(net438),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _2620_ (.A(net438),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _2621_ (.A(net437),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _2622_ (.A(net437),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_2 _2623_ (.A(net443),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_2 _2624_ (.A(net438),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_2 _2625_ (.A(net437),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_2 _2626_ (.A(net443),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _2627_ (.A(net440),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _2628_ (.A(net442),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _2629_ (.A(net440),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _2630_ (.A(net443),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _2631_ (.A(net444),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _2632_ (.A(net442),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _2633_ (.A(net440),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _2634_ (.A(net442),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _2635_ (.A(net442),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _2636_ (.A(net407),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _2637_ (.A(net408),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _2638_ (.A(net407),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _2639_ (.A(net408),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _2640_ (.A(net407),
    .Y(_0178_));
 sky130_fd_sc_hd__nor2_1 _2641_ (.A(\state[4] ),
    .B(\state[0] ),
    .Y(_1922_));
 sky130_fd_sc_hd__and3_2 _2642_ (.A(net264),
    .B(net263),
    .C(_1922_),
    .X(_1923_));
 sky130_fd_sc_hd__clkbuf_2 _2643_ (.A(_1923_),
    .X(_1924_));
 sky130_fd_sc_hd__clkbuf_2 _2644_ (.A(_1924_),
    .X(_1925_));
 sky130_fd_sc_hd__buf_2 _2645_ (.A(_1925_),
    .X(_1926_));
 sky130_fd_sc_hd__nand2_2 _2646_ (.A(net261),
    .B(_1923_),
    .Y(_1927_));
 sky130_fd_sc_hd__buf_2 _2647_ (.A(_1927_),
    .X(_1928_));
 sky130_fd_sc_hd__or2_1 _2648_ (.A(net388),
    .B(net394),
    .X(_1929_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2649_ (.A(_1929_),
    .X(_1930_));
 sky130_fd_sc_hd__clkbuf_2 _2650_ (.A(_1930_),
    .X(_1931_));
 sky130_fd_sc_hd__clkbuf_2 _2651_ (.A(_1931_),
    .X(_1932_));
 sky130_fd_sc_hd__clkbuf_2 _2652_ (.A(_1932_),
    .X(_1933_));
 sky130_fd_sc_hd__clkbuf_2 _2653_ (.A(_1933_),
    .X(_1934_));
 sky130_fd_sc_hd__clkbuf_2 _2654_ (.A(_1934_),
    .X(_1935_));
 sky130_fd_sc_hd__and3_1 _2655_ (.A(net390),
    .B(net396),
    .C(net113),
    .X(_1936_));
 sky130_fd_sc_hd__inv_2 _2656_ (.A(net386),
    .Y(_1937_));
 sky130_fd_sc_hd__clkbuf_2 _2657_ (.A(_1937_),
    .X(_1938_));
 sky130_fd_sc_hd__clkbuf_2 _2658_ (.A(_1938_),
    .X(_1939_));
 sky130_fd_sc_hd__clkbuf_2 _2659_ (.A(_1939_),
    .X(_1940_));
 sky130_fd_sc_hd__clkbuf_2 _2660_ (.A(_1940_),
    .X(_1941_));
 sky130_fd_sc_hd__clkbuf_2 _2661_ (.A(_1941_),
    .X(_1942_));
 sky130_fd_sc_hd__and2b_1 _2662_ (.A_N(net392),
    .B(net386),
    .X(_1943_));
 sky130_fd_sc_hd__clkbuf_2 _2663_ (.A(_1943_),
    .X(_1944_));
 sky130_fd_sc_hd__clkbuf_2 _2664_ (.A(_1944_),
    .X(_1945_));
 sky130_fd_sc_hd__clkbuf_2 _2665_ (.A(_1945_),
    .X(_1946_));
 sky130_fd_sc_hd__nor2_1 _2666_ (.A(net388),
    .B(net394),
    .Y(_1947_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2667_ (.A(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__clkbuf_2 _2668_ (.A(_1948_),
    .X(_1949_));
 sky130_fd_sc_hd__clkbuf_2 _2669_ (.A(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__clkbuf_2 _2670_ (.A(_1950_),
    .X(_1951_));
 sky130_fd_sc_hd__clkbuf_2 _2671_ (.A(_1951_),
    .X(_1952_));
 sky130_fd_sc_hd__a221o_1 _2672_ (.A1(_1942_),
    .A2(net184),
    .B1(_1946_),
    .B2(net149),
    .C1(_1952_),
    .X(_1953_));
 sky130_fd_sc_hd__o22a_2 _2673_ (.A1(net92),
    .A2(_1935_),
    .B1(_1936_),
    .B2(_1953_),
    .X(_1954_));
 sky130_fd_sc_hd__and3_1 _2674_ (.A(net390),
    .B(net396),
    .C(net111),
    .X(_1955_));
 sky130_fd_sc_hd__inv_2 _2675_ (.A(net392),
    .Y(_1956_));
 sky130_fd_sc_hd__buf_2 _2676_ (.A(_1956_),
    .X(_1957_));
 sky130_fd_sc_hd__clkbuf_2 _2677_ (.A(_1957_),
    .X(_1958_));
 sky130_fd_sc_hd__and2b_1 _2678_ (.A_N(net390),
    .B(net396),
    .X(_1959_));
 sky130_fd_sc_hd__a221o_1 _2679_ (.A1(_1958_),
    .A2(net146),
    .B1(net182),
    .B2(_1959_),
    .C1(_1952_),
    .X(_1960_));
 sky130_fd_sc_hd__o22a_1 _2680_ (.A1(net90),
    .A2(_1935_),
    .B1(_1955_),
    .B2(_1960_),
    .X(_1961_));
 sky130_fd_sc_hd__nand2_1 _2681_ (.A(\sum[26] ),
    .B(_1961_),
    .Y(_1962_));
 sky130_fd_sc_hd__and2_1 _2682_ (.A(net386),
    .B(net392),
    .X(_1963_));
 sky130_fd_sc_hd__clkbuf_2 _2683_ (.A(_1963_),
    .X(_1964_));
 sky130_fd_sc_hd__clkbuf_2 _2684_ (.A(_1964_),
    .X(_1965_));
 sky130_fd_sc_hd__clkbuf_2 _2685_ (.A(_1965_),
    .X(_1966_));
 sky130_fd_sc_hd__a221o_1 _2686_ (.A1(_1941_),
    .A2(net179),
    .B1(_1966_),
    .B2(net109),
    .C1(_1951_),
    .X(_1967_));
 sky130_fd_sc_hd__and2_1 _2687_ (.A(net144),
    .B(_1946_),
    .X(_1968_));
 sky130_fd_sc_hd__o22a_1 _2688_ (.A1(net88),
    .A2(_1934_),
    .B1(_1967_),
    .B2(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__nand2_2 _2689_ (.A(\sum[24] ),
    .B(_1969_),
    .Y(_1970_));
 sky130_fd_sc_hd__a22o_1 _2690_ (.A1(_1958_),
    .A2(net143),
    .B1(_1966_),
    .B2(net108),
    .X(_1971_));
 sky130_fd_sc_hd__o21a_1 _2691_ (.A1(_1958_),
    .A2(net178),
    .B1(_1941_),
    .X(_1972_));
 sky130_fd_sc_hd__o22a_1 _2692_ (.A1(net86),
    .A2(_1934_),
    .B1(_1971_),
    .B2(_1972_),
    .X(_1973_));
 sky130_fd_sc_hd__and2_1 _2693_ (.A(\sum[23] ),
    .B(_1973_),
    .X(_1974_));
 sky130_fd_sc_hd__and3_1 _2694_ (.A(net390),
    .B(net396),
    .C(net107),
    .X(_1975_));
 sky130_fd_sc_hd__a221o_1 _2695_ (.A1(_1941_),
    .A2(net177),
    .B1(_1946_),
    .B2(net142),
    .C1(_1951_),
    .X(_1976_));
 sky130_fd_sc_hd__o22a_1 _2696_ (.A1(net85),
    .A2(_1934_),
    .B1(_1975_),
    .B2(_1976_),
    .X(_1977_));
 sky130_fd_sc_hd__nand2_1 _2697_ (.A(\sum[22] ),
    .B(_1977_),
    .Y(_1978_));
 sky130_fd_sc_hd__and3_1 _2698_ (.A(net390),
    .B(net396),
    .C(net106),
    .X(_1979_));
 sky130_fd_sc_hd__a221o_1 _2699_ (.A1(_1941_),
    .A2(net176),
    .B1(_1945_),
    .B2(net141),
    .C1(_1951_),
    .X(_1980_));
 sky130_fd_sc_hd__o22a_1 _2700_ (.A1(net84),
    .A2(_1933_),
    .B1(_1979_),
    .B2(_1980_),
    .X(_1981_));
 sky130_fd_sc_hd__and2_1 _2701_ (.A(\sum[21] ),
    .B(_1981_),
    .X(_1982_));
 sky130_fd_sc_hd__inv_2 _2702_ (.A(_1982_),
    .Y(_1983_));
 sky130_fd_sc_hd__or2_1 _2703_ (.A(net75),
    .B(_1932_),
    .X(_1984_));
 sky130_fd_sc_hd__a22o_1 _2704_ (.A1(_1957_),
    .A2(net132),
    .B1(_1965_),
    .B2(net97),
    .X(_1985_));
 sky130_fd_sc_hd__a211o_1 _2705_ (.A1(_1940_),
    .A2(net167),
    .B1(_1950_),
    .C1(_1985_),
    .X(_1986_));
 sky130_fd_sc_hd__a21oi_1 _2706_ (.A1(_1984_),
    .A2(_1986_),
    .B1(\sum[13] ),
    .Y(_1987_));
 sky130_fd_sc_hd__nand3_1 _2707_ (.A(\sum[13] ),
    .B(_1984_),
    .C(_1986_),
    .Y(_1988_));
 sky130_fd_sc_hd__a22o_1 _2708_ (.A1(_1957_),
    .A2(net131),
    .B1(_1964_),
    .B2(net96),
    .X(_1989_));
 sky130_fd_sc_hd__o21a_1 _2709_ (.A1(_1957_),
    .A2(net166),
    .B1(_1940_),
    .X(_1990_));
 sky130_fd_sc_hd__o22a_1 _2710_ (.A1(net74),
    .A2(_1932_),
    .B1(_1989_),
    .B2(_1990_),
    .X(_1991_));
 sky130_fd_sc_hd__nand2_1 _2711_ (.A(net379),
    .B(_1991_),
    .Y(_1992_));
 sky130_fd_sc_hd__and2_1 _2712_ (.A(_1988_),
    .B(_1992_),
    .X(_1993_));
 sky130_fd_sc_hd__a221o_1 _2713_ (.A1(_1939_),
    .A2(net168),
    .B1(_1964_),
    .B2(net98),
    .C1(_1949_),
    .X(_1994_));
 sky130_fd_sc_hd__a21o_1 _2714_ (.A1(net133),
    .A2(_1944_),
    .B1(_1994_),
    .X(_1995_));
 sky130_fd_sc_hd__or2_1 _2715_ (.A(net77),
    .B(_1932_),
    .X(_1996_));
 sky130_fd_sc_hd__nand3_1 _2716_ (.A(\sum[14] ),
    .B(_1995_),
    .C(_1996_),
    .Y(_1997_));
 sky130_fd_sc_hd__a21o_1 _2717_ (.A1(_1995_),
    .A2(_1996_),
    .B1(\sum[14] ),
    .X(_1998_));
 sky130_fd_sc_hd__nand2_1 _2718_ (.A(_1997_),
    .B(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__a221o_1 _2719_ (.A1(_1938_),
    .A2(net169),
    .B1(_1944_),
    .B2(net134),
    .C1(_1949_),
    .X(_2000_));
 sky130_fd_sc_hd__a21o_1 _2720_ (.A1(net99),
    .A2(_1964_),
    .B1(_2000_),
    .X(_2001_));
 sky130_fd_sc_hd__or2_1 _2721_ (.A(net78),
    .B(_1931_),
    .X(_2002_));
 sky130_fd_sc_hd__a21oi_1 _2722_ (.A1(_2001_),
    .A2(_2002_),
    .B1(\sum[15] ),
    .Y(_2003_));
 sky130_fd_sc_hd__and3_1 _2723_ (.A(\sum[15] ),
    .B(_2001_),
    .C(_2002_),
    .X(_2004_));
 sky130_fd_sc_hd__or2_2 _2724_ (.A(_2003_),
    .B(_2004_),
    .X(_2005_));
 sky130_fd_sc_hd__or2_1 _2725_ (.A(_1999_),
    .B(_2005_),
    .X(_2006_));
 sky130_fd_sc_hd__o21ba_1 _2726_ (.A1(_1997_),
    .A2(_2003_),
    .B1_N(_2004_),
    .X(_2007_));
 sky130_fd_sc_hd__o31a_1 _2727_ (.A1(_1987_),
    .A2(_1993_),
    .A3(_2006_),
    .B1(_2007_),
    .X(_2008_));
 sky130_fd_sc_hd__a221o_1 _2728_ (.A1(_1956_),
    .A2(net129),
    .B1(_1963_),
    .B2(net76),
    .C1(_1949_),
    .X(_2009_));
 sky130_fd_sc_hd__and2_1 _2729_ (.A(_1938_),
    .B(net164),
    .X(_2010_));
 sky130_fd_sc_hd__o22a_1 _2730_ (.A1(net72),
    .A2(_1931_),
    .B1(_2009_),
    .B2(_2010_),
    .X(_2011_));
 sky130_fd_sc_hd__and2_1 _2731_ (.A(\sum[10] ),
    .B(_2011_),
    .X(_2012_));
 sky130_fd_sc_hd__inv_2 _2732_ (.A(_2012_),
    .Y(_2013_));
 sky130_fd_sc_hd__and3_1 _2733_ (.A(net386),
    .B(net392),
    .C(net87),
    .X(_2014_));
 sky130_fd_sc_hd__a221o_1 _2734_ (.A1(_1939_),
    .A2(net165),
    .B1(_1944_),
    .B2(net130),
    .C1(_1949_),
    .X(_2015_));
 sky130_fd_sc_hd__o22a_2 _2735_ (.A1(net73),
    .A2(_1932_),
    .B1(_2014_),
    .B2(_2015_),
    .X(_2016_));
 sky130_fd_sc_hd__nor2_1 _2736_ (.A(net380),
    .B(_2016_),
    .Y(_2017_));
 sky130_fd_sc_hd__nor2_1 _2737_ (.A(\sum[10] ),
    .B(_2011_),
    .Y(_2018_));
 sky130_fd_sc_hd__or2_1 _2738_ (.A(_2012_),
    .B(_2018_),
    .X(_2019_));
 sky130_fd_sc_hd__xnor2_4 _2739_ (.A(net380),
    .B(_2016_),
    .Y(_2020_));
 sky130_fd_sc_hd__or2_1 _2740_ (.A(_2019_),
    .B(_2020_),
    .X(_2021_));
 sky130_fd_sc_hd__and3_1 _2741_ (.A(net389),
    .B(net395),
    .C(net192),
    .X(_2022_));
 sky130_fd_sc_hd__a221o_1 _2742_ (.A1(_1939_),
    .A2(net163),
    .B1(_1944_),
    .B2(net128),
    .C1(_1949_),
    .X(_2023_));
 sky130_fd_sc_hd__o22a_2 _2743_ (.A1(net71),
    .A2(_1932_),
    .B1(_2022_),
    .B2(_2023_),
    .X(_2024_));
 sky130_fd_sc_hd__a22o_1 _2744_ (.A1(_1957_),
    .A2(net127),
    .B1(_1964_),
    .B2(net181),
    .X(_2025_));
 sky130_fd_sc_hd__o21a_1 _2745_ (.A1(_1957_),
    .A2(net162),
    .B1(_1939_),
    .X(_2026_));
 sky130_fd_sc_hd__o22a_1 _2746_ (.A1(net70),
    .A2(_1931_),
    .B1(_2025_),
    .B2(_2026_),
    .X(_2027_));
 sky130_fd_sc_hd__and2_1 _2747_ (.A(\sum[8] ),
    .B(_2027_),
    .X(_2028_));
 sky130_fd_sc_hd__a21o_1 _2748_ (.A1(net382),
    .A2(_2024_),
    .B1(_2028_),
    .X(_2029_));
 sky130_fd_sc_hd__o21ai_1 _2749_ (.A1(net382),
    .A2(_2024_),
    .B1(_2029_),
    .Y(_2030_));
 sky130_fd_sc_hd__nand2_1 _2750_ (.A(net380),
    .B(_2016_),
    .Y(_2031_));
 sky130_fd_sc_hd__o221a_1 _2751_ (.A1(_2013_),
    .A2(_2017_),
    .B1(_2021_),
    .B2(_2030_),
    .C1(_2031_),
    .X(_2032_));
 sky130_fd_sc_hd__and3_1 _2752_ (.A(net386),
    .B(net393),
    .C(net148),
    .X(_2033_));
 sky130_fd_sc_hd__and3b_1 _2753_ (.A_N(net392),
    .B(net123),
    .C(net386),
    .X(_2034_));
 sky130_fd_sc_hd__a2111o_1 _2754_ (.A1(_1937_),
    .A2(net158),
    .B1(_1948_),
    .C1(_2033_),
    .D1(_2034_),
    .X(_2035_));
 sky130_fd_sc_hd__or2_1 _2755_ (.A(net67),
    .B(_1929_),
    .X(_2036_));
 sky130_fd_sc_hd__a21oi_2 _2756_ (.A1(_2035_),
    .A2(_2036_),
    .B1(\sum[5] ),
    .Y(_2037_));
 sky130_fd_sc_hd__a221o_1 _2757_ (.A1(_1956_),
    .A2(net122),
    .B1(_1963_),
    .B2(net137),
    .C1(_1947_),
    .X(_2038_));
 sky130_fd_sc_hd__and2_1 _2758_ (.A(_1937_),
    .B(net157),
    .X(_2039_));
 sky130_fd_sc_hd__o22a_2 _2759_ (.A1(net66),
    .A2(_1930_),
    .B1(_2038_),
    .B2(_2039_),
    .X(_2040_));
 sky130_fd_sc_hd__nand2_1 _2760_ (.A(\sum[4] ),
    .B(_2040_),
    .Y(_2041_));
 sky130_fd_sc_hd__nand3_1 _2761_ (.A(\sum[5] ),
    .B(_2035_),
    .C(_2036_),
    .Y(_2042_));
 sky130_fd_sc_hd__o21a_1 _2762_ (.A1(_2037_),
    .A2(_2041_),
    .B1(_2042_),
    .X(_2043_));
 sky130_fd_sc_hd__and2_1 _2763_ (.A(net124),
    .B(_1943_),
    .X(_2044_));
 sky130_fd_sc_hd__a221o_1 _2764_ (.A1(_1937_),
    .A2(net160),
    .B1(_1963_),
    .B2(net159),
    .C1(_1948_),
    .X(_2045_));
 sky130_fd_sc_hd__o22a_2 _2765_ (.A1(net68),
    .A2(_1930_),
    .B1(_2044_),
    .B2(_2045_),
    .X(_2046_));
 sky130_fd_sc_hd__xnor2_4 _2766_ (.A(net383),
    .B(_2046_),
    .Y(_2047_));
 sky130_fd_sc_hd__and2_1 _2767_ (.A(net161),
    .B(_1959_),
    .X(_2048_));
 sky130_fd_sc_hd__a221o_1 _2768_ (.A1(_1956_),
    .A2(net125),
    .B1(_1963_),
    .B2(net170),
    .C1(_1948_),
    .X(_2049_));
 sky130_fd_sc_hd__o22a_2 _2769_ (.A1(net69),
    .A2(_1930_),
    .B1(_2048_),
    .B2(_2049_),
    .X(_2050_));
 sky130_fd_sc_hd__xnor2_4 _2770_ (.A(\sum[7] ),
    .B(_2050_),
    .Y(_2051_));
 sky130_fd_sc_hd__o211a_1 _2771_ (.A1(\sum[7] ),
    .A2(_2050_),
    .B1(_2046_),
    .C1(net383),
    .X(_2052_));
 sky130_fd_sc_hd__a21oi_1 _2772_ (.A1(\sum[7] ),
    .A2(_2050_),
    .B1(_2052_),
    .Y(_2053_));
 sky130_fd_sc_hd__o31a_1 _2773_ (.A1(_2043_),
    .A2(_2047_),
    .A3(_2051_),
    .B1(_2053_),
    .X(_2054_));
 sky130_fd_sc_hd__a221o_1 _2774_ (.A1(_1938_),
    .A2(net156),
    .B1(_1944_),
    .B2(net121),
    .C1(_1948_),
    .X(_2055_));
 sky130_fd_sc_hd__a21o_1 _2775_ (.A1(net126),
    .A2(_1964_),
    .B1(_2055_),
    .X(_2056_));
 sky130_fd_sc_hd__or2_1 _2776_ (.A(net191),
    .B(_1931_),
    .X(_2057_));
 sky130_fd_sc_hd__a21oi_1 _2777_ (.A1(_2056_),
    .A2(_2057_),
    .B1(\sum[3] ),
    .Y(_2058_));
 sky130_fd_sc_hd__a22o_1 _2778_ (.A1(_1956_),
    .A2(net118),
    .B1(_1963_),
    .B2(net65),
    .X(_2059_));
 sky130_fd_sc_hd__o21a_1 _2779_ (.A1(_1956_),
    .A2(net153),
    .B1(_1938_),
    .X(_2060_));
 sky130_fd_sc_hd__o221a_1 _2780_ (.A1(net188),
    .A2(_1930_),
    .B1(_2059_),
    .B2(_2060_),
    .C1(net385),
    .X(_2061_));
 sky130_fd_sc_hd__or2_1 _2781_ (.A(net189),
    .B(_1929_),
    .X(_2062_));
 sky130_fd_sc_hd__and3b_1 _2782_ (.A_N(net394),
    .B(net119),
    .C(net388),
    .X(_2063_));
 sky130_fd_sc_hd__and3b_1 _2783_ (.A_N(net388),
    .B(net394),
    .C(net154),
    .X(_2064_));
 sky130_fd_sc_hd__and3_1 _2784_ (.A(net388),
    .B(net394),
    .C(net104),
    .X(_2065_));
 sky130_fd_sc_hd__or4_1 _2785_ (.A(_1947_),
    .B(_2063_),
    .C(_2064_),
    .D(_2065_),
    .X(_2066_));
 sky130_fd_sc_hd__a21o_1 _2786_ (.A1(_2062_),
    .A2(_2066_),
    .B1(net384),
    .X(_2067_));
 sky130_fd_sc_hd__and3_1 _2787_ (.A(net384),
    .B(_2062_),
    .C(_2066_),
    .X(_2068_));
 sky130_fd_sc_hd__a21oi_2 _2788_ (.A1(_2061_),
    .A2(_2067_),
    .B1(_2068_),
    .Y(_2069_));
 sky130_fd_sc_hd__and3_1 _2789_ (.A(net387),
    .B(net393),
    .C(net115),
    .X(_2070_));
 sky130_fd_sc_hd__and3b_1 _2790_ (.A_N(net392),
    .B(net120),
    .C(net387),
    .X(_2071_));
 sky130_fd_sc_hd__a2111o_1 _2791_ (.A1(_1938_),
    .A2(net155),
    .B1(_1948_),
    .C1(_2070_),
    .D1(_2071_),
    .X(_2072_));
 sky130_fd_sc_hd__or2_1 _2792_ (.A(net190),
    .B(_1930_),
    .X(_2073_));
 sky130_fd_sc_hd__nand3_1 _2793_ (.A(\sum[2] ),
    .B(_2072_),
    .C(_2073_),
    .Y(_2074_));
 sky130_fd_sc_hd__a21o_1 _2794_ (.A1(_2072_),
    .A2(_2073_),
    .B1(\sum[2] ),
    .X(_2075_));
 sky130_fd_sc_hd__nand2_1 _2795_ (.A(_2074_),
    .B(_2075_),
    .Y(_2076_));
 sky130_fd_sc_hd__nand3_1 _2796_ (.A(\sum[3] ),
    .B(_2056_),
    .C(_2057_),
    .Y(_2077_));
 sky130_fd_sc_hd__o211a_1 _2797_ (.A1(_2069_),
    .A2(_2076_),
    .B1(_2077_),
    .C1(_2074_),
    .X(_2078_));
 sky130_fd_sc_hd__xnor2_4 _2798_ (.A(\sum[4] ),
    .B(_2040_),
    .Y(_2079_));
 sky130_fd_sc_hd__or2b_1 _2799_ (.A(_2037_),
    .B_N(_2042_),
    .X(_2080_));
 sky130_fd_sc_hd__or4_1 _2800_ (.A(_2079_),
    .B(_2080_),
    .C(_2047_),
    .D(_2051_),
    .X(_2081_));
 sky130_fd_sc_hd__or3_2 _2801_ (.A(_2058_),
    .B(_2078_),
    .C(_2081_),
    .X(_2082_));
 sky130_fd_sc_hd__nor2_1 _2802_ (.A(\sum[8] ),
    .B(_2027_),
    .Y(_2083_));
 sky130_fd_sc_hd__or2_1 _2803_ (.A(_2028_),
    .B(_2083_),
    .X(_2084_));
 sky130_fd_sc_hd__xnor2_2 _2804_ (.A(\sum[9] ),
    .B(_2024_),
    .Y(_2085_));
 sky130_fd_sc_hd__a2111o_1 _2805_ (.A1(_2054_),
    .A2(_2082_),
    .B1(_2084_),
    .C1(_2085_),
    .D1(_2021_),
    .X(_2086_));
 sky130_fd_sc_hd__and3_1 _2806_ (.A(_2008_),
    .B(_2032_),
    .C(_2086_),
    .X(_2087_));
 sky130_fd_sc_hd__or2b_1 _2807_ (.A(_1987_),
    .B_N(_1988_),
    .X(_2088_));
 sky130_fd_sc_hd__or2_1 _2808_ (.A(\sum[12] ),
    .B(_1991_),
    .X(_2089_));
 sky130_fd_sc_hd__nand2_1 _2809_ (.A(_1992_),
    .B(_2089_),
    .Y(_2090_));
 sky130_fd_sc_hd__o31a_1 _2810_ (.A1(_2006_),
    .A2(_2088_),
    .A3(_2090_),
    .B1(_2008_),
    .X(_2091_));
 sky130_fd_sc_hd__and3_1 _2811_ (.A(net390),
    .B(net396),
    .C(net100),
    .X(_2092_));
 sky130_fd_sc_hd__a221o_1 _2812_ (.A1(_1940_),
    .A2(net171),
    .B1(_1945_),
    .B2(net135),
    .C1(_1950_),
    .X(_2093_));
 sky130_fd_sc_hd__o22a_1 _2813_ (.A1(net79),
    .A2(_1933_),
    .B1(_2092_),
    .B2(_2093_),
    .X(_2094_));
 sky130_fd_sc_hd__nand2_1 _2814_ (.A(\sum[16] ),
    .B(_2094_),
    .Y(_2095_));
 sky130_fd_sc_hd__or2_1 _2815_ (.A(\sum[16] ),
    .B(_2094_),
    .X(_2096_));
 sky130_fd_sc_hd__nand2_2 _2816_ (.A(_2095_),
    .B(_2096_),
    .Y(_2097_));
 sky130_fd_sc_hd__a221o_1 _2817_ (.A1(_1939_),
    .A2(net172),
    .B1(_1945_),
    .B2(net136),
    .C1(_1950_),
    .X(_2098_));
 sky130_fd_sc_hd__a21o_1 _2818_ (.A1(net101),
    .A2(_1965_),
    .B1(_2098_),
    .X(_2099_));
 sky130_fd_sc_hd__or2_1 _2819_ (.A(net80),
    .B(_1933_),
    .X(_2100_));
 sky130_fd_sc_hd__and3_1 _2820_ (.A(\sum[17] ),
    .B(_2099_),
    .C(_2100_),
    .X(_2101_));
 sky130_fd_sc_hd__a21oi_2 _2821_ (.A1(_2099_),
    .A2(_2100_),
    .B1(\sum[17] ),
    .Y(_2102_));
 sky130_fd_sc_hd__or2_1 _2822_ (.A(_2101_),
    .B(_2102_),
    .X(_2103_));
 sky130_fd_sc_hd__and2_1 _2823_ (.A(net138),
    .B(_1945_),
    .X(_2104_));
 sky130_fd_sc_hd__a221o_1 _2824_ (.A1(_1940_),
    .A2(net173),
    .B1(_1965_),
    .B2(net102),
    .C1(_1950_),
    .X(_2105_));
 sky130_fd_sc_hd__o22a_1 _2825_ (.A1(net81),
    .A2(_1933_),
    .B1(_2104_),
    .B2(_2105_),
    .X(_2106_));
 sky130_fd_sc_hd__nand2_1 _2826_ (.A(\sum[18] ),
    .B(_2106_),
    .Y(_2107_));
 sky130_fd_sc_hd__or2_1 _2827_ (.A(\sum[18] ),
    .B(_2106_),
    .X(_2108_));
 sky130_fd_sc_hd__nand2_2 _2828_ (.A(_2107_),
    .B(_2108_),
    .Y(_2109_));
 sky130_fd_sc_hd__and2_1 _2829_ (.A(net139),
    .B(_1945_),
    .X(_2110_));
 sky130_fd_sc_hd__a221o_1 _2830_ (.A1(_1940_),
    .A2(net174),
    .B1(_1965_),
    .B2(net103),
    .C1(_1950_),
    .X(_2111_));
 sky130_fd_sc_hd__o22a_2 _2831_ (.A1(net82),
    .A2(_1933_),
    .B1(_2110_),
    .B2(_2111_),
    .X(_2112_));
 sky130_fd_sc_hd__xnor2_4 _2832_ (.A(net378),
    .B(_2112_),
    .Y(_2113_));
 sky130_fd_sc_hd__or4_1 _2833_ (.A(_2097_),
    .B(_2103_),
    .C(_2109_),
    .D(_2113_),
    .X(_2114_));
 sky130_fd_sc_hd__or3_1 _2834_ (.A(_2087_),
    .B(_2091_),
    .C(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__nor2_1 _2835_ (.A(_2109_),
    .B(_2113_),
    .Y(_2116_));
 sky130_fd_sc_hd__o21bai_1 _2836_ (.A1(_2095_),
    .A2(_2102_),
    .B1_N(_2101_),
    .Y(_2117_));
 sky130_fd_sc_hd__o211a_1 _2837_ (.A1(\sum[19] ),
    .A2(_2112_),
    .B1(_2106_),
    .C1(\sum[18] ),
    .X(_2118_));
 sky130_fd_sc_hd__a221oi_2 _2838_ (.A1(net378),
    .A2(_2112_),
    .B1(_2116_),
    .B2(_2117_),
    .C1(_2118_),
    .Y(_2119_));
 sky130_fd_sc_hd__nor2_1 _2839_ (.A(\sum[21] ),
    .B(_1981_),
    .Y(_2120_));
 sky130_fd_sc_hd__or2_2 _2840_ (.A(_1982_),
    .B(_2120_),
    .X(_2121_));
 sky130_fd_sc_hd__a221o_1 _2841_ (.A1(_1958_),
    .A2(net140),
    .B1(_1965_),
    .B2(net105),
    .C1(_1951_),
    .X(_2122_));
 sky130_fd_sc_hd__a21o_1 _2842_ (.A1(_1941_),
    .A2(net175),
    .B1(_2122_),
    .X(_2123_));
 sky130_fd_sc_hd__o21a_1 _2843_ (.A1(net83),
    .A2(_1934_),
    .B1(_2123_),
    .X(_2124_));
 sky130_fd_sc_hd__and2_1 _2844_ (.A(\sum[20] ),
    .B(_2124_),
    .X(_2125_));
 sky130_fd_sc_hd__nor2_1 _2845_ (.A(\sum[20] ),
    .B(_2124_),
    .Y(_2126_));
 sky130_fd_sc_hd__or2_1 _2846_ (.A(_2125_),
    .B(_2126_),
    .X(_2127_));
 sky130_fd_sc_hd__a211o_1 _2847_ (.A1(_2115_),
    .A2(_2119_),
    .B1(_2121_),
    .C1(_2127_),
    .X(_2128_));
 sky130_fd_sc_hd__or2b_1 _2848_ (.A(_2120_),
    .B_N(_2125_),
    .X(_2129_));
 sky130_fd_sc_hd__or2_1 _2849_ (.A(\sum[22] ),
    .B(_1977_),
    .X(_2130_));
 sky130_fd_sc_hd__nand2_2 _2850_ (.A(_1978_),
    .B(_2130_),
    .Y(_2131_));
 sky130_fd_sc_hd__a31o_1 _2851_ (.A1(_1983_),
    .A2(_2128_),
    .A3(_2129_),
    .B1(_2131_),
    .X(_2132_));
 sky130_fd_sc_hd__nor2_1 _2852_ (.A(\sum[23] ),
    .B(_1973_),
    .Y(_2133_));
 sky130_fd_sc_hd__or2_1 _2853_ (.A(_1974_),
    .B(_2133_),
    .X(_2134_));
 sky130_fd_sc_hd__a21oi_1 _2854_ (.A1(_1978_),
    .A2(_2132_),
    .B1(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hd__or2_1 _2855_ (.A(\sum[24] ),
    .B(_1969_),
    .X(_2136_));
 sky130_fd_sc_hd__nand2_1 _2856_ (.A(_1970_),
    .B(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__o21bai_2 _2857_ (.A1(_1974_),
    .A2(_2135_),
    .B1_N(_2137_),
    .Y(_2138_));
 sky130_fd_sc_hd__a221o_1 _2858_ (.A1(_1942_),
    .A2(net180),
    .B1(_1946_),
    .B2(net145),
    .C1(_1951_),
    .X(_2139_));
 sky130_fd_sc_hd__a21o_1 _2859_ (.A1(net110),
    .A2(_1966_),
    .B1(_2139_),
    .X(_2140_));
 sky130_fd_sc_hd__or2_1 _2860_ (.A(net89),
    .B(_1934_),
    .X(_2141_));
 sky130_fd_sc_hd__nand3_1 _2861_ (.A(\sum[25] ),
    .B(_2140_),
    .C(_2141_),
    .Y(_2142_));
 sky130_fd_sc_hd__a21oi_1 _2862_ (.A1(_2140_),
    .A2(_2141_),
    .B1(\sum[25] ),
    .Y(_2143_));
 sky130_fd_sc_hd__or2_1 _2863_ (.A(\sum[26] ),
    .B(_1961_),
    .X(_2144_));
 sky130_fd_sc_hd__nand2_2 _2864_ (.A(_1962_),
    .B(_2144_),
    .Y(_2145_));
 sky130_fd_sc_hd__a311o_1 _2865_ (.A1(_1970_),
    .A2(_2138_),
    .A3(_2142_),
    .B1(_2143_),
    .C1(_2145_),
    .X(_2146_));
 sky130_fd_sc_hd__a221o_1 _2866_ (.A1(_1958_),
    .A2(net147),
    .B1(_1966_),
    .B2(net112),
    .C1(_1952_),
    .X(_2147_));
 sky130_fd_sc_hd__and2_1 _2867_ (.A(_1942_),
    .B(net183),
    .X(_2148_));
 sky130_fd_sc_hd__o22a_1 _2868_ (.A1(net91),
    .A2(_1935_),
    .B1(_2147_),
    .B2(_2148_),
    .X(_2149_));
 sky130_fd_sc_hd__nand2_1 _2869_ (.A(\sum[27] ),
    .B(_2149_),
    .Y(_2150_));
 sky130_fd_sc_hd__xnor2_4 _2870_ (.A(\sum[28] ),
    .B(_1954_),
    .Y(_2151_));
 sky130_fd_sc_hd__nor2_1 _2871_ (.A(\sum[27] ),
    .B(_2149_),
    .Y(_2152_));
 sky130_fd_sc_hd__a311o_1 _2872_ (.A1(_1962_),
    .A2(_2146_),
    .A3(_2150_),
    .B1(_2151_),
    .C1(_2152_),
    .X(_2153_));
 sky130_fd_sc_hd__a21bo_2 _2873_ (.A1(\sum[28] ),
    .A2(_1954_),
    .B1_N(_2153_),
    .X(_2154_));
 sky130_fd_sc_hd__or2_1 _2874_ (.A(net93),
    .B(_1935_),
    .X(_2155_));
 sky130_fd_sc_hd__a221o_1 _2875_ (.A1(_1958_),
    .A2(net150),
    .B1(_1966_),
    .B2(net114),
    .C1(_1952_),
    .X(_2156_));
 sky130_fd_sc_hd__a21o_1 _2876_ (.A1(_1942_),
    .A2(net185),
    .B1(_2156_),
    .X(_2157_));
 sky130_fd_sc_hd__a21oi_2 _2877_ (.A1(_2155_),
    .A2(_2157_),
    .B1(\sum[29] ),
    .Y(_2158_));
 sky130_fd_sc_hd__and3_1 _2878_ (.A(\sum[29] ),
    .B(_2155_),
    .C(_2157_),
    .X(_2159_));
 sky130_fd_sc_hd__nor2_2 _2879_ (.A(_2158_),
    .B(_2159_),
    .Y(_2160_));
 sky130_fd_sc_hd__xnor2_4 _2880_ (.A(_2154_),
    .B(_2160_),
    .Y(_2161_));
 sky130_fd_sc_hd__or2_1 _2881_ (.A(net325),
    .B(net332),
    .X(_2162_));
 sky130_fd_sc_hd__xor2_1 _2882_ (.A(\workunit1[31] ),
    .B(net337),
    .X(_2163_));
 sky130_fd_sc_hd__nand2_1 _2883_ (.A(net328),
    .B(_2163_),
    .Y(_2164_));
 sky130_fd_sc_hd__or2_1 _2884_ (.A(net328),
    .B(_2163_),
    .X(_2165_));
 sky130_fd_sc_hd__nand2_1 _2885_ (.A(_2164_),
    .B(_2165_),
    .Y(_2166_));
 sky130_fd_sc_hd__xor2_1 _2886_ (.A(net324),
    .B(net340),
    .X(_2167_));
 sky130_fd_sc_hd__nand2_1 _2887_ (.A(net332),
    .B(_2167_),
    .Y(_2168_));
 sky130_fd_sc_hd__or2_1 _2888_ (.A(net332),
    .B(net350),
    .X(_2169_));
 sky130_fd_sc_hd__nand2_1 _2889_ (.A(net332),
    .B(net350),
    .Y(_2170_));
 sky130_fd_sc_hd__a21o_1 _2890_ (.A1(_2169_),
    .A2(_2170_),
    .B1(net342),
    .X(_2171_));
 sky130_fd_sc_hd__or2_1 _2891_ (.A(net334),
    .B(net352),
    .X(_2172_));
 sky130_fd_sc_hd__nand2_1 _2892_ (.A(net334),
    .B(net352),
    .Y(_2173_));
 sky130_fd_sc_hd__a21o_1 _2893_ (.A1(_2172_),
    .A2(_2173_),
    .B1(net344),
    .X(_2174_));
 sky130_fd_sc_hd__nand3_1 _2894_ (.A(net342),
    .B(_2169_),
    .C(_2170_),
    .Y(_2175_));
 sky130_fd_sc_hd__a21boi_1 _2895_ (.A1(_2171_),
    .A2(_2174_),
    .B1_N(_2175_),
    .Y(_2176_));
 sky130_fd_sc_hd__xor2_1 _2896_ (.A(net346),
    .B(net364),
    .X(_2177_));
 sky130_fd_sc_hd__or2_1 _2897_ (.A(net344),
    .B(net362),
    .X(_2178_));
 sky130_fd_sc_hd__nand2_1 _2898_ (.A(net344),
    .B(net362),
    .Y(_2179_));
 sky130_fd_sc_hd__a21o_1 _2899_ (.A1(_2178_),
    .A2(_2179_),
    .B1(net354),
    .X(_2180_));
 sky130_fd_sc_hd__and3_1 _2900_ (.A(net355),
    .B(_2178_),
    .C(_2179_),
    .X(_2181_));
 sky130_fd_sc_hd__a31oi_2 _2901_ (.A1(net356),
    .A2(_2177_),
    .A3(_2180_),
    .B1(_2181_),
    .Y(_2182_));
 sky130_fd_sc_hd__or2_1 _2902_ (.A(net354),
    .B(net372),
    .X(_2183_));
 sky130_fd_sc_hd__nand2_1 _2903_ (.A(net354),
    .B(net372),
    .Y(_2184_));
 sky130_fd_sc_hd__and3_1 _2904_ (.A(net365),
    .B(_2183_),
    .C(_2184_),
    .X(_2185_));
 sky130_fd_sc_hd__a21oi_1 _2905_ (.A1(_2183_),
    .A2(_2184_),
    .B1(net365),
    .Y(_2186_));
 sky130_fd_sc_hd__or2_1 _2906_ (.A(_2185_),
    .B(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__or2_1 _2907_ (.A(net352),
    .B(net371),
    .X(_2188_));
 sky130_fd_sc_hd__nand2_1 _2908_ (.A(net352),
    .B(net370),
    .Y(_2189_));
 sky130_fd_sc_hd__a21o_1 _2909_ (.A1(_2188_),
    .A2(_2189_),
    .B1(net362),
    .X(_0353_));
 sky130_fd_sc_hd__nand3_1 _2910_ (.A(net363),
    .B(_2188_),
    .C(_2189_),
    .Y(_0354_));
 sky130_fd_sc_hd__nand2_1 _2911_ (.A(_0353_),
    .B(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__xor2_1 _2912_ (.A(net350),
    .B(net369),
    .X(_0356_));
 sky130_fd_sc_hd__nand2_1 _2913_ (.A(net360),
    .B(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__or2_1 _2914_ (.A(net360),
    .B(_0356_),
    .X(_0358_));
 sky130_fd_sc_hd__nand2_1 _2915_ (.A(_0357_),
    .B(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__or2_1 _2916_ (.A(net348),
    .B(net366),
    .X(_0360_));
 sky130_fd_sc_hd__nand2_1 _2917_ (.A(net348),
    .B(net366),
    .Y(_0361_));
 sky130_fd_sc_hd__and3_1 _2918_ (.A(net359),
    .B(_0360_),
    .C(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__a21oi_1 _2919_ (.A1(_0360_),
    .A2(_0361_),
    .B1(net358),
    .Y(_0363_));
 sky130_fd_sc_hd__or2_1 _2920_ (.A(_0362_),
    .B(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__nor2_1 _2921_ (.A(_0359_),
    .B(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__or2_1 _2922_ (.A(net356),
    .B(net373),
    .X(_0366_));
 sky130_fd_sc_hd__nand2_1 _2923_ (.A(net356),
    .B(net373),
    .Y(_0367_));
 sky130_fd_sc_hd__a21o_1 _2924_ (.A1(_0366_),
    .A2(_0367_),
    .B1(net367),
    .X(_0368_));
 sky130_fd_sc_hd__or2_1 _2925_ (.A(net359),
    .B(net374),
    .X(_0369_));
 sky130_fd_sc_hd__nand2_1 _2926_ (.A(net358),
    .B(net374),
    .Y(_0370_));
 sky130_fd_sc_hd__a21o_1 _2927_ (.A1(_0369_),
    .A2(_0370_),
    .B1(net368),
    .X(_0371_));
 sky130_fd_sc_hd__or2_1 _2928_ (.A(net360),
    .B(net375),
    .X(_0372_));
 sky130_fd_sc_hd__nand2_1 _2929_ (.A(net360),
    .B(net375),
    .Y(_0373_));
 sky130_fd_sc_hd__a21o_1 _2930_ (.A1(_0372_),
    .A2(_0373_),
    .B1(net370),
    .X(_0374_));
 sky130_fd_sc_hd__or2_1 _2931_ (.A(net364),
    .B(\workunit1[3] ),
    .X(_0375_));
 sky130_fd_sc_hd__xor2_1 _2932_ (.A(net369),
    .B(net375),
    .X(_0376_));
 sky130_fd_sc_hd__and2_1 _2933_ (.A(net369),
    .B(net375),
    .X(_0377_));
 sky130_fd_sc_hd__a31o_1 _2934_ (.A1(net370),
    .A2(net377),
    .A3(_0376_),
    .B1(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__or2_1 _2935_ (.A(net367),
    .B(\workunit1[2] ),
    .X(_0379_));
 sky130_fd_sc_hd__nand2_1 _2936_ (.A(net367),
    .B(\workunit1[2] ),
    .Y(_0380_));
 sky130_fd_sc_hd__a21bo_1 _2937_ (.A1(_0378_),
    .A2(_0379_),
    .B1_N(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__nand2_1 _2938_ (.A(net365),
    .B(\workunit1[3] ),
    .Y(_0382_));
 sky130_fd_sc_hd__a21bo_1 _2939_ (.A1(_0375_),
    .A2(_0381_),
    .B1_N(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__or2_1 _2940_ (.A(net363),
    .B(net376),
    .X(_0384_));
 sky130_fd_sc_hd__nand2_1 _2941_ (.A(net363),
    .B(net377),
    .Y(_0385_));
 sky130_fd_sc_hd__and3_1 _2942_ (.A(\workunit1[4] ),
    .B(_0384_),
    .C(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__a21oi_1 _2943_ (.A1(_0384_),
    .A2(_0385_),
    .B1(\workunit1[4] ),
    .Y(_0387_));
 sky130_fd_sc_hd__or2_1 _2944_ (.A(_0386_),
    .B(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__inv_2 _2945_ (.A(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__nand3_1 _2946_ (.A(net370),
    .B(_0372_),
    .C(_0373_),
    .Y(_0390_));
 sky130_fd_sc_hd__inv_2 _2947_ (.A(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__a211o_1 _2948_ (.A1(_0383_),
    .A2(_0389_),
    .B1(_0391_),
    .C1(_0386_),
    .X(_0392_));
 sky130_fd_sc_hd__and3_1 _2949_ (.A(net368),
    .B(_0369_),
    .C(_0370_),
    .X(_0393_));
 sky130_fd_sc_hd__a31o_1 _2950_ (.A1(_0371_),
    .A2(_0374_),
    .A3(_0392_),
    .B1(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__and3_1 _2951_ (.A(net367),
    .B(_0366_),
    .C(_0367_),
    .X(_0395_));
 sky130_fd_sc_hd__a21o_1 _2952_ (.A1(_0368_),
    .A2(_0394_),
    .B1(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__or4bb_1 _2953_ (.A(_2187_),
    .B(_0355_),
    .C_N(_0365_),
    .D_N(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__or2b_1 _2954_ (.A(_2185_),
    .B_N(_0354_),
    .X(_0398_));
 sky130_fd_sc_hd__a31o_1 _2955_ (.A1(_0353_),
    .A2(_0365_),
    .A3(_0398_),
    .B1(_0362_),
    .X(_0399_));
 sky130_fd_sc_hd__o21ba_1 _2956_ (.A1(_0357_),
    .A2(_0363_),
    .B1_N(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__nand2_1 _2957_ (.A(net357),
    .B(_2177_),
    .Y(_0401_));
 sky130_fd_sc_hd__or2_1 _2958_ (.A(net357),
    .B(_2177_),
    .X(_0402_));
 sky130_fd_sc_hd__nand2_1 _2959_ (.A(_0401_),
    .B(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__or2b_1 _2960_ (.A(_2181_),
    .B_N(_2180_),
    .X(_0404_));
 sky130_fd_sc_hd__a211o_1 _2961_ (.A1(_0397_),
    .A2(_0400_),
    .B1(_0403_),
    .C1(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__or2_1 _2962_ (.A(net339),
    .B(net359),
    .X(_0406_));
 sky130_fd_sc_hd__nand2_1 _2963_ (.A(net339),
    .B(net359),
    .Y(_0407_));
 sky130_fd_sc_hd__a21oi_1 _2964_ (.A1(_0406_),
    .A2(_0407_),
    .B1(net350),
    .Y(_0408_));
 sky130_fd_sc_hd__xor2_1 _2965_ (.A(net341),
    .B(net361),
    .X(_0409_));
 sky130_fd_sc_hd__nand2_1 _2966_ (.A(net353),
    .B(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__nand3_1 _2967_ (.A(net351),
    .B(_0406_),
    .C(_0407_),
    .Y(_0411_));
 sky130_fd_sc_hd__o21a_1 _2968_ (.A1(_0408_),
    .A2(_0410_),
    .B1(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__nor2_1 _2969_ (.A(net352),
    .B(_0409_),
    .Y(_0413_));
 sky130_fd_sc_hd__o21a_1 _2970_ (.A1(_0408_),
    .A2(_0413_),
    .B1(_0411_),
    .X(_0414_));
 sky130_fd_sc_hd__a31o_1 _2971_ (.A1(_2182_),
    .A2(_0405_),
    .A3(_0412_),
    .B1(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__xor2_1 _2972_ (.A(net338),
    .B(net356),
    .X(_0416_));
 sky130_fd_sc_hd__and2_1 _2973_ (.A(net348),
    .B(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__nor2_1 _2974_ (.A(net348),
    .B(_0416_),
    .Y(_0418_));
 sky130_fd_sc_hd__or2_1 _2975_ (.A(_0417_),
    .B(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__or2_1 _2976_ (.A(net336),
    .B(net354),
    .X(_0420_));
 sky130_fd_sc_hd__nand2_1 _2977_ (.A(net336),
    .B(net354),
    .Y(_0421_));
 sky130_fd_sc_hd__a21oi_1 _2978_ (.A1(_0420_),
    .A2(_0421_),
    .B1(net346),
    .Y(_0422_));
 sky130_fd_sc_hd__nand3_1 _2979_ (.A(net346),
    .B(_0420_),
    .C(_0421_),
    .Y(_0423_));
 sky130_fd_sc_hd__or2b_1 _2980_ (.A(_0422_),
    .B_N(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__or2_1 _2981_ (.A(_0419_),
    .B(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__inv_2 _2982_ (.A(_0417_),
    .Y(_0426_));
 sky130_fd_sc_hd__a21o_1 _2983_ (.A1(_0426_),
    .A2(_0423_),
    .B1(_0422_),
    .X(_0427_));
 sky130_fd_sc_hd__nand3_1 _2984_ (.A(net344),
    .B(_2172_),
    .C(_2173_),
    .Y(_0428_));
 sky130_fd_sc_hd__and2_1 _2985_ (.A(_2175_),
    .B(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__o211a_1 _2986_ (.A1(_0415_),
    .A2(_0425_),
    .B1(_0427_),
    .C1(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__xor2_1 _2987_ (.A(net330),
    .B(net349),
    .X(_0431_));
 sky130_fd_sc_hd__nand2_1 _2988_ (.A(net339),
    .B(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__or2_1 _2989_ (.A(net339),
    .B(_0431_),
    .X(_0433_));
 sky130_fd_sc_hd__nand2_1 _2990_ (.A(_0432_),
    .B(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__or2_1 _2991_ (.A(net328),
    .B(net346),
    .X(_0435_));
 sky130_fd_sc_hd__nand2_1 _2992_ (.A(net328),
    .B(net347),
    .Y(_0436_));
 sky130_fd_sc_hd__nand3_1 _2993_ (.A(net338),
    .B(_0435_),
    .C(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__a21o_1 _2994_ (.A1(_0435_),
    .A2(_0436_),
    .B1(net338),
    .X(_0438_));
 sky130_fd_sc_hd__nand2_1 _2995_ (.A(_0437_),
    .B(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__a21bo_1 _2996_ (.A1(_0432_),
    .A2(_0437_),
    .B1_N(_0438_),
    .X(_0440_));
 sky130_fd_sc_hd__o41a_2 _2997_ (.A1(_2176_),
    .A2(_0430_),
    .A3(_0434_),
    .A4(_0439_),
    .B1(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__or2_1 _2998_ (.A(net325),
    .B(net342),
    .X(_0442_));
 sky130_fd_sc_hd__nand2_1 _2999_ (.A(net325),
    .B(net341),
    .Y(_0443_));
 sky130_fd_sc_hd__nand3_2 _3000_ (.A(net335),
    .B(_0442_),
    .C(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__or2_1 _3001_ (.A(net327),
    .B(net345),
    .X(_0445_));
 sky130_fd_sc_hd__nand2_1 _3002_ (.A(net327),
    .B(net345),
    .Y(_0446_));
 sky130_fd_sc_hd__and3_1 _3003_ (.A(net336),
    .B(_0445_),
    .C(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__inv_2 _3004_ (.A(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__a21oi_1 _3005_ (.A1(_0442_),
    .A2(_0443_),
    .B1(net334),
    .Y(_0449_));
 sky130_fd_sc_hd__a21o_1 _3006_ (.A1(_0444_),
    .A2(_0448_),
    .B1(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__a21oi_1 _3007_ (.A1(_0445_),
    .A2(_0446_),
    .B1(net336),
    .Y(_0451_));
 sky130_fd_sc_hd__or2_1 _3008_ (.A(_0449_),
    .B(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__or2_1 _3009_ (.A(net332),
    .B(_2167_),
    .X(_0453_));
 sky130_fd_sc_hd__nand2_1 _3010_ (.A(_2168_),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__a221o_1 _3011_ (.A1(_0441_),
    .A2(_0450_),
    .B1(_0452_),
    .B2(_0444_),
    .C1(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__or2_1 _3012_ (.A(net323),
    .B(net338),
    .X(_0456_));
 sky130_fd_sc_hd__nand2_1 _3013_ (.A(net323),
    .B(\workunit1[21] ),
    .Y(_0457_));
 sky130_fd_sc_hd__nand3_1 _3014_ (.A(net330),
    .B(_0456_),
    .C(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__a21oi_1 _3015_ (.A1(_0456_),
    .A2(_0457_),
    .B1(net330),
    .Y(_0459_));
 sky130_fd_sc_hd__a31o_1 _3016_ (.A1(_2168_),
    .A2(_0455_),
    .A3(_0458_),
    .B1(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__o21ai_1 _3017_ (.A1(_2166_),
    .A2(_0460_),
    .B1(_2164_),
    .Y(_0461_));
 sky130_fd_sc_hd__or2_1 _3018_ (.A(net327),
    .B(net335),
    .X(_0462_));
 sky130_fd_sc_hd__and2_1 _3019_ (.A(net326),
    .B(net335),
    .X(_0463_));
 sky130_fd_sc_hd__a21o_1 _3020_ (.A1(_0461_),
    .A2(_0462_),
    .B1(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__nand2_1 _3021_ (.A(\workunit1[28] ),
    .B(net332),
    .Y(_0465_));
 sky130_fd_sc_hd__a21boi_1 _3022_ (.A1(_2162_),
    .A2(_0464_),
    .B1_N(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__nor2_1 _3023_ (.A(net324),
    .B(net330),
    .Y(_0467_));
 sky130_fd_sc_hd__nand2_1 _3024_ (.A(net324),
    .B(net330),
    .Y(_0468_));
 sky130_fd_sc_hd__and2b_1 _3025_ (.A_N(_0467_),
    .B(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__xnor2_1 _3026_ (.A(_0466_),
    .B(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__xnor2_1 _3027_ (.A(_2161_),
    .B(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__inv_2 _3028_ (.A(_2143_),
    .Y(_0472_));
 sky130_fd_sc_hd__nand2_1 _3029_ (.A(_2142_),
    .B(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__nand3_2 _3030_ (.A(_1970_),
    .B(_2138_),
    .C(_0473_),
    .Y(_0474_));
 sky130_fd_sc_hd__a21o_1 _3031_ (.A1(_1970_),
    .A2(_2138_),
    .B1(_0473_),
    .X(_0475_));
 sky130_fd_sc_hd__nand2_1 _3032_ (.A(_0474_),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__nand2_1 _3033_ (.A(_2168_),
    .B(_0455_),
    .Y(_0477_));
 sky130_fd_sc_hd__and3_1 _3034_ (.A(net330),
    .B(_0456_),
    .C(_0457_),
    .X(_0478_));
 sky130_fd_sc_hd__nor2_1 _3035_ (.A(_0478_),
    .B(_0459_),
    .Y(_0479_));
 sky130_fd_sc_hd__xor2_1 _3036_ (.A(_0477_),
    .B(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__xnor2_2 _3037_ (.A(_0476_),
    .B(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__or2_1 _3038_ (.A(_2176_),
    .B(_0430_),
    .X(_0482_));
 sky130_fd_sc_hd__o21a_1 _3039_ (.A1(_0482_),
    .A2(_0434_),
    .B1(_0432_),
    .X(_0483_));
 sky130_fd_sc_hd__a21oi_1 _3040_ (.A1(_2115_),
    .A2(_2119_),
    .B1(_2127_),
    .Y(_0484_));
 sky130_fd_sc_hd__nor2_2 _3041_ (.A(_2125_),
    .B(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__xnor2_4 _3042_ (.A(_2121_),
    .B(_0485_),
    .Y(_0486_));
 sky130_fd_sc_hd__xnor2_1 _3043_ (.A(_0439_),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__xor2_1 _3044_ (.A(_0483_),
    .B(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__nand2_1 _3045_ (.A(_2171_),
    .B(_2175_),
    .Y(_0489_));
 sky130_fd_sc_hd__o21ai_1 _3046_ (.A1(_0415_),
    .A2(_0425_),
    .B1(_0427_),
    .Y(_0490_));
 sky130_fd_sc_hd__a21bo_1 _3047_ (.A1(_2174_),
    .A2(_0490_),
    .B1_N(_0428_),
    .X(_0491_));
 sky130_fd_sc_hd__xor2_2 _3048_ (.A(_0489_),
    .B(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__o31a_2 _3049_ (.A1(_2097_),
    .A2(_2087_),
    .A3(_2091_),
    .B1(_2095_),
    .X(_0493_));
 sky130_fd_sc_hd__o21bai_4 _3050_ (.A1(_2102_),
    .A2(_0493_),
    .B1_N(_2101_),
    .Y(_0494_));
 sky130_fd_sc_hd__a21bo_1 _3051_ (.A1(_2108_),
    .A2(_0494_),
    .B1_N(_2107_),
    .X(_0495_));
 sky130_fd_sc_hd__xor2_4 _3052_ (.A(_2113_),
    .B(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__xnor2_2 _3053_ (.A(_0492_),
    .B(_0496_),
    .Y(_0497_));
 sky130_fd_sc_hd__a21o_1 _3054_ (.A1(_2032_),
    .A2(_2086_),
    .B1(_2090_),
    .X(_0498_));
 sky130_fd_sc_hd__a21oi_2 _3055_ (.A1(_1993_),
    .A2(_0498_),
    .B1(_1987_),
    .Y(_0499_));
 sky130_fd_sc_hd__a21bo_1 _3056_ (.A1(_1998_),
    .A2(_0499_),
    .B1_N(_1997_),
    .X(_0500_));
 sky130_fd_sc_hd__xor2_4 _3057_ (.A(_2005_),
    .B(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__inv_2 _3058_ (.A(_0411_),
    .Y(_0502_));
 sky130_fd_sc_hd__nor2_1 _3059_ (.A(_0502_),
    .B(_0408_),
    .Y(_0503_));
 sky130_fd_sc_hd__or2_1 _3060_ (.A(net352),
    .B(_0409_),
    .X(_0504_));
 sky130_fd_sc_hd__nand2_1 _3061_ (.A(_0410_),
    .B(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__a21o_1 _3062_ (.A1(_2182_),
    .A2(_0405_),
    .B1(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__nand3_1 _3063_ (.A(_0410_),
    .B(_0503_),
    .C(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__a21o_1 _3064_ (.A1(_0410_),
    .A2(_0506_),
    .B1(_0503_),
    .X(_0508_));
 sky130_fd_sc_hd__and3_1 _3065_ (.A(_0501_),
    .B(_0507_),
    .C(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__a21oi_1 _3066_ (.A1(_0507_),
    .A2(_0508_),
    .B1(_0501_),
    .Y(_0510_));
 sky130_fd_sc_hd__inv_2 _3067_ (.A(\state[3] ),
    .Y(_0511_));
 sky130_fd_sc_hd__and2_1 _3068_ (.A(net264),
    .B(_1922_),
    .X(_0512_));
 sky130_fd_sc_hd__nand2_4 _3069_ (.A(net263),
    .B(_0512_),
    .Y(_0513_));
 sky130_fd_sc_hd__nor2_1 _3070_ (.A(_0511_),
    .B(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__buf_1 _3071_ (.A(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__inv_2 _3072_ (.A(_0353_),
    .Y(_0516_));
 sky130_fd_sc_hd__inv_2 _3073_ (.A(_2187_),
    .Y(_0517_));
 sky130_fd_sc_hd__a21oi_1 _3074_ (.A1(_0396_),
    .A2(_0517_),
    .B1(_0398_),
    .Y(_0518_));
 sky130_fd_sc_hd__or2_1 _3075_ (.A(_0516_),
    .B(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__xnor2_1 _3076_ (.A(_0359_),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__a211o_1 _3077_ (.A1(_2054_),
    .A2(_2082_),
    .B1(_2084_),
    .C1(_2085_),
    .X(_0521_));
 sky130_fd_sc_hd__a21oi_1 _3078_ (.A1(_0521_),
    .A2(_2030_),
    .B1(_2019_),
    .Y(_0522_));
 sky130_fd_sc_hd__and3_1 _3079_ (.A(_0521_),
    .B(_2030_),
    .C(_2019_),
    .X(_0523_));
 sky130_fd_sc_hd__or2_2 _3080_ (.A(_0522_),
    .B(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__xnor2_2 _3081_ (.A(_0520_),
    .B(_0524_),
    .Y(_0525_));
 sky130_fd_sc_hd__a21oi_1 _3082_ (.A1(_2054_),
    .A2(_2082_),
    .B1(_2084_),
    .Y(_0526_));
 sky130_fd_sc_hd__nor2_1 _3083_ (.A(_2028_),
    .B(_0526_),
    .Y(_0527_));
 sky130_fd_sc_hd__xnor2_2 _3084_ (.A(_2085_),
    .B(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__a21oi_1 _3085_ (.A1(_0396_),
    .A2(_0517_),
    .B1(_2185_),
    .Y(_0529_));
 sky130_fd_sc_hd__xnor2_1 _3086_ (.A(_0355_),
    .B(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__xnor2_1 _3087_ (.A(_0528_),
    .B(_0530_),
    .Y(_0531_));
 sky130_fd_sc_hd__xnor2_2 _3088_ (.A(_0383_),
    .B(_0388_),
    .Y(_0532_));
 sky130_fd_sc_hd__or2_2 _3089_ (.A(_2058_),
    .B(_2078_),
    .X(_0533_));
 sky130_fd_sc_hd__xnor2_4 _3090_ (.A(_2079_),
    .B(_0533_),
    .Y(_0534_));
 sky130_fd_sc_hd__xnor2_4 _3091_ (.A(_0532_),
    .B(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__a21o_1 _3092_ (.A1(_0383_),
    .A2(_0389_),
    .B1(_0386_),
    .X(_0536_));
 sky130_fd_sc_hd__nand2_1 _3093_ (.A(_0390_),
    .B(_0374_),
    .Y(_0537_));
 sky130_fd_sc_hd__xnor2_1 _3094_ (.A(_0536_),
    .B(_0537_),
    .Y(_0538_));
 sky130_fd_sc_hd__o31a_1 _3095_ (.A1(_2079_),
    .A2(_2058_),
    .A3(_2078_),
    .B1(_2041_),
    .X(_0539_));
 sky130_fd_sc_hd__xnor2_2 _3096_ (.A(_2080_),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__xnor2_1 _3097_ (.A(_0538_),
    .B(_0540_),
    .Y(_0541_));
 sky130_fd_sc_hd__nand2_1 _3098_ (.A(_0382_),
    .B(_0375_),
    .Y(_0542_));
 sky130_fd_sc_hd__xnor2_1 _3099_ (.A(_0542_),
    .B(_0381_),
    .Y(_0543_));
 sky130_fd_sc_hd__o21a_1 _3100_ (.A1(_2069_),
    .A2(_2076_),
    .B1(_2074_),
    .X(_0544_));
 sky130_fd_sc_hd__a21o_1 _3101_ (.A1(_2056_),
    .A2(_2057_),
    .B1(\sum[3] ),
    .X(_0545_));
 sky130_fd_sc_hd__nand2_1 _3102_ (.A(_2077_),
    .B(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__xnor2_2 _3103_ (.A(_0544_),
    .B(_0546_),
    .Y(_0547_));
 sky130_fd_sc_hd__xnor2_2 _3104_ (.A(_0543_),
    .B(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__nand2_1 _3105_ (.A(net370),
    .B(net376),
    .Y(_0549_));
 sky130_fd_sc_hd__or2_1 _3106_ (.A(net370),
    .B(net376),
    .X(_0550_));
 sky130_fd_sc_hd__nand2_2 _3107_ (.A(_0549_),
    .B(_0550_),
    .Y(_0551_));
 sky130_fd_sc_hd__o22a_2 _3108_ (.A1(net188),
    .A2(_1931_),
    .B1(_2059_),
    .B2(_2060_),
    .X(_0552_));
 sky130_fd_sc_hd__xnor2_4 _3109_ (.A(net385),
    .B(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__xor2_4 _3110_ (.A(_0551_),
    .B(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__and2_1 _3111_ (.A(_1927_),
    .B(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__a21oi_1 _3112_ (.A1(_2062_),
    .A2(_2066_),
    .B1(net384),
    .Y(_0556_));
 sky130_fd_sc_hd__or3b_2 _3113_ (.A(_2068_),
    .B(_0556_),
    .C_N(_2061_),
    .X(_0557_));
 sky130_fd_sc_hd__xnor2_1 _3114_ (.A(_0549_),
    .B(_0376_),
    .Y(_0558_));
 sky130_fd_sc_hd__o21bai_2 _3115_ (.A1(_2068_),
    .A2(_0556_),
    .B1_N(_2061_),
    .Y(_0559_));
 sky130_fd_sc_hd__and3_1 _3116_ (.A(_0557_),
    .B(_0558_),
    .C(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__a21oi_2 _3117_ (.A1(_0557_),
    .A2(_0559_),
    .B1(_0558_),
    .Y(_0561_));
 sky130_fd_sc_hd__nor2_1 _3118_ (.A(_0560_),
    .B(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__nand2_1 _3119_ (.A(_0380_),
    .B(_0379_),
    .Y(_0563_));
 sky130_fd_sc_hd__xor2_1 _3120_ (.A(_0378_),
    .B(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__xor2_2 _3121_ (.A(_2069_),
    .B(_2076_),
    .X(_0565_));
 sky130_fd_sc_hd__xnor2_2 _3122_ (.A(_0564_),
    .B(_0565_),
    .Y(_0566_));
 sky130_fd_sc_hd__o31a_1 _3123_ (.A1(_0555_),
    .A2(_0562_),
    .A3(_0566_),
    .B1(_1927_),
    .X(_0567_));
 sky130_fd_sc_hd__a21o_1 _3124_ (.A1(_1928_),
    .A2(_0548_),
    .B1(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__a211oi_2 _3125_ (.A1(_1928_),
    .A2(_0535_),
    .B1(_0541_),
    .C1(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__or2b_1 _3126_ (.A(_0393_),
    .B_N(_0371_),
    .X(_0570_));
 sky130_fd_sc_hd__nand2_1 _3127_ (.A(_0374_),
    .B(_0392_),
    .Y(_0571_));
 sky130_fd_sc_hd__xnor2_1 _3128_ (.A(_0570_),
    .B(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__o311a_1 _3129_ (.A1(_2079_),
    .A2(_2058_),
    .A3(_2078_),
    .B1(_2042_),
    .C1(_2041_),
    .X(_0573_));
 sky130_fd_sc_hd__nor2_2 _3130_ (.A(_2037_),
    .B(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__xor2_4 _3131_ (.A(_0574_),
    .B(_2047_),
    .X(_0575_));
 sky130_fd_sc_hd__xnor2_2 _3132_ (.A(_0572_),
    .B(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__and2b_1 _3133_ (.A_N(_0395_),
    .B(_0368_),
    .X(_0577_));
 sky130_fd_sc_hd__xnor2_1 _3134_ (.A(_0577_),
    .B(_0394_),
    .Y(_0578_));
 sky130_fd_sc_hd__nand2_1 _3135_ (.A(net383),
    .B(_2046_),
    .Y(_0579_));
 sky130_fd_sc_hd__o31a_2 _3136_ (.A1(_2037_),
    .A2(_0573_),
    .A3(_2047_),
    .B1(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__xnor2_4 _3137_ (.A(_2051_),
    .B(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__xnor2_2 _3138_ (.A(_0578_),
    .B(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__a31o_1 _3139_ (.A1(_0569_),
    .A2(_0576_),
    .A3(_0582_),
    .B1(_0514_),
    .X(_0583_));
 sky130_fd_sc_hd__xnor2_1 _3140_ (.A(_0396_),
    .B(_0517_),
    .Y(_0584_));
 sky130_fd_sc_hd__and3_1 _3141_ (.A(_2054_),
    .B(_2082_),
    .C(_2084_),
    .X(_0585_));
 sky130_fd_sc_hd__or2_1 _3142_ (.A(_0526_),
    .B(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__xnor2_1 _3143_ (.A(_0584_),
    .B(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__or2_1 _3144_ (.A(_0515_),
    .B(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__o211a_1 _3145_ (.A1(_0515_),
    .A2(_0531_),
    .B1(_0583_),
    .C1(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__nor2_2 _3146_ (.A(_2012_),
    .B(_0522_),
    .Y(_0590_));
 sky130_fd_sc_hd__xnor2_4 _3147_ (.A(_2020_),
    .B(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__o31a_1 _3148_ (.A1(_0516_),
    .A2(_0359_),
    .A3(_0518_),
    .B1(_0357_),
    .X(_0592_));
 sky130_fd_sc_hd__xnor2_1 _3149_ (.A(_0364_),
    .B(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__xnor2_1 _3150_ (.A(_0591_),
    .B(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__o211a_1 _3151_ (.A1(_0515_),
    .A2(_0525_),
    .B1(_0589_),
    .C1(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__a21o_1 _3152_ (.A1(_0397_),
    .A2(_0400_),
    .B1(_0403_),
    .X(_0596_));
 sky130_fd_sc_hd__nand3_1 _3153_ (.A(_0401_),
    .B(_0596_),
    .C(_0404_),
    .Y(_0597_));
 sky130_fd_sc_hd__a21o_1 _3154_ (.A1(_0401_),
    .A2(_0596_),
    .B1(_0404_),
    .X(_0598_));
 sky130_fd_sc_hd__nand2_1 _3155_ (.A(_1992_),
    .B(_0498_),
    .Y(_0599_));
 sky130_fd_sc_hd__xor2_2 _3156_ (.A(_2088_),
    .B(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__a21o_1 _3157_ (.A1(_0597_),
    .A2(_0598_),
    .B1(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__nand3_1 _3158_ (.A(_0600_),
    .B(_0597_),
    .C(_0598_),
    .Y(_0602_));
 sky130_fd_sc_hd__nand3_1 _3159_ (.A(_0397_),
    .B(_0400_),
    .C(_0403_),
    .Y(_0603_));
 sky130_fd_sc_hd__nand2_1 _3160_ (.A(_0596_),
    .B(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__nand3_1 _3161_ (.A(_2032_),
    .B(_2086_),
    .C(_2090_),
    .Y(_0605_));
 sky130_fd_sc_hd__nand2_2 _3162_ (.A(_0498_),
    .B(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__xnor2_1 _3163_ (.A(_0604_),
    .B(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__and3_1 _3164_ (.A(_0601_),
    .B(_0602_),
    .C(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__nand3_1 _3165_ (.A(_2182_),
    .B(_0405_),
    .C(_0505_),
    .Y(_0609_));
 sky130_fd_sc_hd__nand2_1 _3166_ (.A(_0506_),
    .B(_0609_),
    .Y(_0610_));
 sky130_fd_sc_hd__xnor2_2 _3167_ (.A(_1999_),
    .B(_0499_),
    .Y(_0611_));
 sky130_fd_sc_hd__xor2_1 _3168_ (.A(_0610_),
    .B(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__o2111a_1 _3169_ (.A1(_0509_),
    .A2(_0510_),
    .B1(_0595_),
    .C1(_0608_),
    .D1(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__xnor2_1 _3170_ (.A(_0415_),
    .B(_0419_),
    .Y(_0614_));
 sky130_fd_sc_hd__nor2_2 _3171_ (.A(_2087_),
    .B(_2091_),
    .Y(_0615_));
 sky130_fd_sc_hd__xor2_4 _3172_ (.A(_2097_),
    .B(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__xnor2_2 _3173_ (.A(_0614_),
    .B(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__o21ai_1 _3174_ (.A1(_0415_),
    .A2(_0419_),
    .B1(_0426_),
    .Y(_0618_));
 sky130_fd_sc_hd__xnor2_2 _3175_ (.A(_2103_),
    .B(_0493_),
    .Y(_0619_));
 sky130_fd_sc_hd__xor2_1 _3176_ (.A(_0424_),
    .B(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__xnor2_1 _3177_ (.A(_0618_),
    .B(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__nand2_1 _3178_ (.A(_2174_),
    .B(_0428_),
    .Y(_0622_));
 sky130_fd_sc_hd__xnor2_1 _3179_ (.A(_0490_),
    .B(_0622_),
    .Y(_0623_));
 sky130_fd_sc_hd__xnor2_4 _3180_ (.A(_2109_),
    .B(_0494_),
    .Y(_0624_));
 sky130_fd_sc_hd__xnor2_1 _3181_ (.A(_0623_),
    .B(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__and4_1 _3182_ (.A(_0613_),
    .B(_0617_),
    .C(_0621_),
    .D(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__xnor2_1 _3183_ (.A(_0482_),
    .B(_0434_),
    .Y(_0627_));
 sky130_fd_sc_hd__and3_1 _3184_ (.A(_2115_),
    .B(_2119_),
    .C(_2127_),
    .X(_0628_));
 sky130_fd_sc_hd__or2_2 _3185_ (.A(_0484_),
    .B(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__xnor2_1 _3186_ (.A(_0627_),
    .B(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__and4b_1 _3187_ (.A_N(_0488_),
    .B(_0497_),
    .C(_0626_),
    .D(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__or2_1 _3188_ (.A(_0447_),
    .B(_0451_),
    .X(_0632_));
 sky130_fd_sc_hd__xnor2_1 _3189_ (.A(_0441_),
    .B(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__nand3_2 _3190_ (.A(_1983_),
    .B(_2128_),
    .C(_2129_),
    .Y(_0634_));
 sky130_fd_sc_hd__xor2_4 _3191_ (.A(_2131_),
    .B(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__xnor2_2 _3192_ (.A(_0633_),
    .B(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__o21ai_1 _3193_ (.A1(_0441_),
    .A2(_0451_),
    .B1(_0448_),
    .Y(_0637_));
 sky130_fd_sc_hd__inv_2 _3194_ (.A(_0444_),
    .Y(_0638_));
 sky130_fd_sc_hd__nor2_1 _3195_ (.A(_0638_),
    .B(_0449_),
    .Y(_0639_));
 sky130_fd_sc_hd__and3_1 _3196_ (.A(_2134_),
    .B(_1978_),
    .C(_2132_),
    .X(_0640_));
 sky130_fd_sc_hd__or2_2 _3197_ (.A(_2135_),
    .B(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__xnor2_1 _3198_ (.A(_0639_),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__xnor2_2 _3199_ (.A(_0637_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__a22o_1 _3200_ (.A1(_0441_),
    .A2(_0450_),
    .B1(_0452_),
    .B2(_0444_),
    .X(_0644_));
 sky130_fd_sc_hd__xor2_1 _3201_ (.A(_0454_),
    .B(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__or3b_1 _3202_ (.A(_1974_),
    .B(_2135_),
    .C_N(_2137_),
    .X(_0646_));
 sky130_fd_sc_hd__and2_2 _3203_ (.A(_2138_),
    .B(_0646_),
    .X(_0647_));
 sky130_fd_sc_hd__xnor2_1 _3204_ (.A(_0645_),
    .B(_0647_),
    .Y(_0648_));
 sky130_fd_sc_hd__nand4_1 _3205_ (.A(_0631_),
    .B(_0636_),
    .C(_0643_),
    .D(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__xor2_2 _3206_ (.A(_2166_),
    .B(_0460_),
    .X(_0650_));
 sky130_fd_sc_hd__a31o_1 _3207_ (.A1(_1970_),
    .A2(_2138_),
    .A3(_2142_),
    .B1(_2143_),
    .X(_0651_));
 sky130_fd_sc_hd__xnor2_4 _3208_ (.A(_2145_),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__xnor2_2 _3209_ (.A(_0650_),
    .B(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__o31a_1 _3210_ (.A1(_0481_),
    .A2(_0649_),
    .A3(_0653_),
    .B1(_1928_),
    .X(_0654_));
 sky130_fd_sc_hd__nand2_2 _3211_ (.A(_1962_),
    .B(_2146_),
    .Y(_0655_));
 sky130_fd_sc_hd__and2b_1 _3212_ (.A_N(_2152_),
    .B(_2150_),
    .X(_0656_));
 sky130_fd_sc_hd__xnor2_4 _3213_ (.A(_0655_),
    .B(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__or2b_1 _3214_ (.A(_0463_),
    .B_N(_0462_),
    .X(_0658_));
 sky130_fd_sc_hd__xnor2_1 _3215_ (.A(_0461_),
    .B(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__xnor2_2 _3216_ (.A(_0657_),
    .B(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__nor2_1 _3217_ (.A(_0654_),
    .B(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__nand2_1 _3218_ (.A(_0465_),
    .B(_2162_),
    .Y(_0662_));
 sky130_fd_sc_hd__xor2_1 _3219_ (.A(_0662_),
    .B(_0464_),
    .X(_0663_));
 sky130_fd_sc_hd__a31o_1 _3220_ (.A1(_1962_),
    .A2(_2146_),
    .A3(_2150_),
    .B1(_2152_),
    .X(_0664_));
 sky130_fd_sc_hd__xnor2_4 _3221_ (.A(_2151_),
    .B(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__xnor2_1 _3222_ (.A(_0663_),
    .B(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3223_ (.A(_0515_),
    .X(_0667_));
 sky130_fd_sc_hd__clkbuf_2 _3224_ (.A(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__clkbuf_2 _3225_ (.A(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__a21o_1 _3226_ (.A1(_0661_),
    .A2(_0666_),
    .B1(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__a21bo_1 _3227_ (.A1(_1928_),
    .A2(_0471_),
    .B1_N(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__nand2_1 _3228_ (.A(net323),
    .B(net328),
    .Y(_0672_));
 sky130_fd_sc_hd__or2_1 _3229_ (.A(\workunit1[30] ),
    .B(net328),
    .X(_0673_));
 sky130_fd_sc_hd__nand2_1 _3230_ (.A(_0672_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__o21ai_1 _3231_ (.A1(_0466_),
    .A2(_0467_),
    .B1(_0468_),
    .Y(_0675_));
 sky130_fd_sc_hd__xnor2_1 _3232_ (.A(_0674_),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__and3_1 _3233_ (.A(net391),
    .B(net397),
    .C(net116),
    .X(_0677_));
 sky130_fd_sc_hd__a221o_1 _3234_ (.A1(_1942_),
    .A2(net186),
    .B1(_1946_),
    .B2(net151),
    .C1(_1952_),
    .X(_0678_));
 sky130_fd_sc_hd__o22a_1 _3235_ (.A1(net94),
    .A2(_1935_),
    .B1(_0677_),
    .B2(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__nand2_1 _3236_ (.A(\sum[30] ),
    .B(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__or2_1 _3237_ (.A(\sum[30] ),
    .B(_0679_),
    .X(_0681_));
 sky130_fd_sc_hd__nand2_2 _3238_ (.A(_0680_),
    .B(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__nor2_1 _3239_ (.A(_2154_),
    .B(_2159_),
    .Y(_0683_));
 sky130_fd_sc_hd__nor2_2 _3240_ (.A(_2158_),
    .B(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__xnor2_4 _3241_ (.A(_0682_),
    .B(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__xnor2_1 _3242_ (.A(_0676_),
    .B(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__xnor2_1 _3243_ (.A(_0671_),
    .B(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__nand2_1 _3244_ (.A(\workunit2[30] ),
    .B(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__or2_1 _3245_ (.A(net266),
    .B(_0687_),
    .X(_0689_));
 sky130_fd_sc_hd__nand2_1 _3246_ (.A(_0688_),
    .B(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__or2_1 _3247_ (.A(_0669_),
    .B(_0661_),
    .X(_0691_));
 sky130_fd_sc_hd__xnor2_1 _3248_ (.A(_0691_),
    .B(_0666_),
    .Y(_0692_));
 sky130_fd_sc_hd__or2b_1 _3249_ (.A(_0692_),
    .B_N(\workunit2[28] ),
    .X(_0693_));
 sky130_fd_sc_hd__a21oi_1 _3250_ (.A1(_0631_),
    .A2(_0636_),
    .B1(_0668_),
    .Y(_0694_));
 sky130_fd_sc_hd__xnor2_2 _3251_ (.A(_0643_),
    .B(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__xnor2_1 _3252_ (.A(net279),
    .B(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__nor2_1 _3253_ (.A(_0668_),
    .B(_0631_),
    .Y(_0697_));
 sky130_fd_sc_hd__xnor2_2 _3254_ (.A(_0636_),
    .B(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__xnor2_2 _3255_ (.A(net281),
    .B(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__nor2_1 _3256_ (.A(_0696_),
    .B(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__clkbuf_2 _3257_ (.A(_0667_),
    .X(_0701_));
 sky130_fd_sc_hd__a21o_1 _3258_ (.A1(_0497_),
    .A2(_0626_),
    .B1(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__xnor2_1 _3259_ (.A(_0630_),
    .B(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__and2b_1 _3260_ (.A_N(_0703_),
    .B(net284),
    .X(_0704_));
 sky130_fd_sc_hd__a31o_1 _3261_ (.A1(_0497_),
    .A2(_0626_),
    .A3(_0630_),
    .B1(_0701_),
    .X(_0705_));
 sky130_fd_sc_hd__xnor2_1 _3262_ (.A(_0488_),
    .B(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__nand2_1 _3263_ (.A(net282),
    .B(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__inv_2 _3264_ (.A(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__nor2_1 _3265_ (.A(net283),
    .B(_0706_),
    .Y(_0709_));
 sky130_fd_sc_hd__o21ba_1 _3266_ (.A1(_0704_),
    .A2(_0708_),
    .B1_N(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__and2b_1 _3267_ (.A_N(net285),
    .B(_0703_),
    .X(_0711_));
 sky130_fd_sc_hd__nor2_1 _3268_ (.A(_0704_),
    .B(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__and2b_1 _3269_ (.A_N(_0709_),
    .B(_0707_),
    .X(_0713_));
 sky130_fd_sc_hd__and4bb_1 _3270_ (.A_N(_0696_),
    .B_N(_0699_),
    .C(_0712_),
    .D(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__nor2_1 _3271_ (.A(_0701_),
    .B(_0626_),
    .Y(_0715_));
 sky130_fd_sc_hd__xnor2_2 _3272_ (.A(_0497_),
    .B(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__xnor2_1 _3273_ (.A(net287),
    .B(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__a31o_1 _3274_ (.A1(_0613_),
    .A2(_0617_),
    .A3(_0621_),
    .B1(_0667_),
    .X(_0718_));
 sky130_fd_sc_hd__xor2_1 _3275_ (.A(_0625_),
    .B(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__nand2_1 _3276_ (.A(net290),
    .B(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__or2_1 _3277_ (.A(net289),
    .B(_0719_),
    .X(_0721_));
 sky130_fd_sc_hd__nand2_1 _3278_ (.A(_0720_),
    .B(_0721_),
    .Y(_0722_));
 sky130_fd_sc_hd__or2_1 _3279_ (.A(_0717_),
    .B(_0722_),
    .X(_0723_));
 sky130_fd_sc_hd__a21o_1 _3280_ (.A1(_0613_),
    .A2(_0617_),
    .B1(_0668_),
    .X(_0724_));
 sky130_fd_sc_hd__xor2_1 _3281_ (.A(_0621_),
    .B(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__nor2_1 _3282_ (.A(net291),
    .B(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__and2_1 _3283_ (.A(net291),
    .B(_0725_),
    .X(_0727_));
 sky130_fd_sc_hd__nor2_1 _3284_ (.A(_0668_),
    .B(_0613_),
    .Y(_0728_));
 sky130_fd_sc_hd__xnor2_1 _3285_ (.A(_0617_),
    .B(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__and2_1 _3286_ (.A(net293),
    .B(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__nor2_1 _3287_ (.A(_0727_),
    .B(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__o21ba_1 _3288_ (.A1(net287),
    .A2(_0716_),
    .B1_N(_0720_),
    .X(_0732_));
 sky130_fd_sc_hd__a21oi_1 _3289_ (.A1(net287),
    .A2(_0716_),
    .B1(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__o31ai_4 _3290_ (.A1(_0723_),
    .A2(_0726_),
    .A3(_0731_),
    .B1(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__o211a_1 _3291_ (.A1(net279),
    .A2(_0695_),
    .B1(_0698_),
    .C1(net281),
    .X(_0735_));
 sky130_fd_sc_hd__a21o_1 _3292_ (.A1(\workunit2[23] ),
    .A2(_0695_),
    .B1(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__a221oi_2 _3293_ (.A1(_0700_),
    .A2(_0710_),
    .B1(_0714_),
    .B2(_0734_),
    .C1(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__nor2_1 _3294_ (.A(_0509_),
    .B(_0510_),
    .Y(_0738_));
 sky130_fd_sc_hd__and2_1 _3295_ (.A(_0595_),
    .B(_0608_),
    .X(_0739_));
 sky130_fd_sc_hd__a21o_1 _3296_ (.A1(_0739_),
    .A2(_0612_),
    .B1(_0701_),
    .X(_0740_));
 sky130_fd_sc_hd__xnor2_1 _3297_ (.A(_0738_),
    .B(_0740_),
    .Y(_0741_));
 sky130_fd_sc_hd__and2_1 _3298_ (.A(net295),
    .B(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__nor2_1 _3299_ (.A(_0667_),
    .B(_0739_),
    .Y(_0743_));
 sky130_fd_sc_hd__xnor2_1 _3300_ (.A(_0612_),
    .B(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__nand2_1 _3301_ (.A(net297),
    .B(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__nand2_1 _3302_ (.A(_0601_),
    .B(_0602_),
    .Y(_0746_));
 sky130_fd_sc_hd__a21o_1 _3303_ (.A1(_0595_),
    .A2(_0607_),
    .B1(_0701_),
    .X(_0747_));
 sky130_fd_sc_hd__xnor2_1 _3304_ (.A(_0746_),
    .B(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__nand2_1 _3305_ (.A(net299),
    .B(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__or2_1 _3306_ (.A(_0667_),
    .B(_0595_),
    .X(_0750_));
 sky130_fd_sc_hd__xor2_1 _3307_ (.A(_0607_),
    .B(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__nand2_1 _3308_ (.A(net301),
    .B(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__o21ai_1 _3309_ (.A1(_0667_),
    .A2(_0525_),
    .B1(_0589_),
    .Y(_0753_));
 sky130_fd_sc_hd__xnor2_1 _3310_ (.A(_0753_),
    .B(_0594_),
    .Y(_0754_));
 sky130_fd_sc_hd__nand2_1 _3311_ (.A(net304),
    .B(_0754_),
    .Y(_0755_));
 sky130_fd_sc_hd__xor2_1 _3312_ (.A(_0525_),
    .B(_0589_),
    .X(_0756_));
 sky130_fd_sc_hd__nand2_1 _3313_ (.A(net305),
    .B(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__nand2_1 _3314_ (.A(_0583_),
    .B(_0588_),
    .Y(_0758_));
 sky130_fd_sc_hd__xnor2_1 _3315_ (.A(_0531_),
    .B(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__nand2_1 _3316_ (.A(net307),
    .B(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__xor2_1 _3317_ (.A(_0587_),
    .B(_0583_),
    .X(_0761_));
 sky130_fd_sc_hd__nand2_1 _3318_ (.A(net309),
    .B(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__a21oi_1 _3319_ (.A1(_0569_),
    .A2(_0576_),
    .B1(_0515_),
    .Y(_0763_));
 sky130_fd_sc_hd__xnor2_1 _3320_ (.A(_0763_),
    .B(_0582_),
    .Y(_0764_));
 sky130_fd_sc_hd__and2_1 _3321_ (.A(net312),
    .B(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__nor2_1 _3322_ (.A(_0515_),
    .B(_0569_),
    .Y(_0766_));
 sky130_fd_sc_hd__xnor2_2 _3323_ (.A(_0576_),
    .B(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__nand2_1 _3324_ (.A(net314),
    .B(_0767_),
    .Y(_0768_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3325_ (.A(_0511_),
    .X(_0769_));
 sky130_fd_sc_hd__o221a_1 _3326_ (.A1(_0769_),
    .A2(_0513_),
    .B1(_0568_),
    .B2(_0535_),
    .C1(_0541_),
    .X(_0770_));
 sky130_fd_sc_hd__nor2_1 _3327_ (.A(_0569_),
    .B(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__and2_1 _3328_ (.A(net316),
    .B(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__xor2_2 _3329_ (.A(_0568_),
    .B(_0535_),
    .X(_0773_));
 sky130_fd_sc_hd__nand2_1 _3330_ (.A(net317),
    .B(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__xor2_2 _3331_ (.A(_0567_),
    .B(_0548_),
    .X(_0775_));
 sky130_fd_sc_hd__nand2_1 _3332_ (.A(net318),
    .B(_0775_),
    .Y(_0776_));
 sky130_fd_sc_hd__a211o_1 _3333_ (.A1(_1927_),
    .A2(_0562_),
    .B1(_0566_),
    .C1(_0555_),
    .X(_0777_));
 sky130_fd_sc_hd__o211ai_2 _3334_ (.A1(_0554_),
    .A2(_0562_),
    .B1(_0566_),
    .C1(_1928_),
    .Y(_0778_));
 sky130_fd_sc_hd__nand3_1 _3335_ (.A(net319),
    .B(_0777_),
    .C(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__and3_1 _3336_ (.A(net319),
    .B(_0777_),
    .C(_0778_),
    .X(_0780_));
 sky130_fd_sc_hd__nand2_1 _3337_ (.A(\workunit2[0] ),
    .B(_0554_),
    .Y(_0781_));
 sky130_fd_sc_hd__inv_2 _3338_ (.A(net321),
    .Y(_0782_));
 sky130_fd_sc_hd__o211ai_2 _3339_ (.A1(_0560_),
    .A2(_0561_),
    .B1(_1927_),
    .C1(_0554_),
    .Y(_0783_));
 sky130_fd_sc_hd__a211o_1 _3340_ (.A1(_1927_),
    .A2(_0554_),
    .B1(_0560_),
    .C1(_0561_),
    .X(_0784_));
 sky130_fd_sc_hd__and3_1 _3341_ (.A(_0782_),
    .B(_0783_),
    .C(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__a21oi_1 _3342_ (.A1(_0783_),
    .A2(_0784_),
    .B1(_0782_),
    .Y(_0786_));
 sky130_fd_sc_hd__o21ba_1 _3343_ (.A1(_0781_),
    .A2(_0785_),
    .B1_N(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__a21oi_1 _3344_ (.A1(_0777_),
    .A2(_0778_),
    .B1(net319),
    .Y(_0788_));
 sky130_fd_sc_hd__or3_1 _3345_ (.A(_0780_),
    .B(_0787_),
    .C(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__xnor2_1 _3346_ (.A(net318),
    .B(_0775_),
    .Y(_0790_));
 sky130_fd_sc_hd__a21o_1 _3347_ (.A1(_0779_),
    .A2(_0789_),
    .B1(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__xnor2_1 _3348_ (.A(net317),
    .B(_0773_),
    .Y(_0792_));
 sky130_fd_sc_hd__a21o_1 _3349_ (.A1(_0776_),
    .A2(_0791_),
    .B1(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__xnor2_1 _3350_ (.A(net316),
    .B(_0771_),
    .Y(_0794_));
 sky130_fd_sc_hd__a21oi_1 _3351_ (.A1(_0774_),
    .A2(_0793_),
    .B1(_0794_),
    .Y(_0795_));
 sky130_fd_sc_hd__xnor2_1 _3352_ (.A(net314),
    .B(_0767_),
    .Y(_0796_));
 sky130_fd_sc_hd__o21bai_1 _3353_ (.A1(_0772_),
    .A2(_0795_),
    .B1_N(_0796_),
    .Y(_0797_));
 sky130_fd_sc_hd__nor2_1 _3354_ (.A(net312),
    .B(_0764_),
    .Y(_0798_));
 sky130_fd_sc_hd__or2_1 _3355_ (.A(_0765_),
    .B(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__a21oi_1 _3356_ (.A1(_0768_),
    .A2(_0797_),
    .B1(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__or2_1 _3357_ (.A(net310),
    .B(_0761_),
    .X(_0801_));
 sky130_fd_sc_hd__and2_1 _3358_ (.A(_0762_),
    .B(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__o21ai_2 _3359_ (.A1(_0765_),
    .A2(_0800_),
    .B1(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__nor2_1 _3360_ (.A(net307),
    .B(_0759_),
    .Y(_0804_));
 sky130_fd_sc_hd__or2_1 _3361_ (.A(net305),
    .B(_0756_),
    .X(_0805_));
 sky130_fd_sc_hd__and2_1 _3362_ (.A(_0757_),
    .B(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__inv_2 _3363_ (.A(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__a311o_1 _3364_ (.A1(_0760_),
    .A2(_0762_),
    .A3(_0803_),
    .B1(_0804_),
    .C1(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__nor2_1 _3365_ (.A(net304),
    .B(_0754_),
    .Y(_0809_));
 sky130_fd_sc_hd__xnor2_1 _3366_ (.A(net301),
    .B(_0751_),
    .Y(_0810_));
 sky130_fd_sc_hd__a311o_1 _3367_ (.A1(_0755_),
    .A2(_0757_),
    .A3(_0808_),
    .B1(_0809_),
    .C1(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__nor2_1 _3368_ (.A(net299),
    .B(_0748_),
    .Y(_0812_));
 sky130_fd_sc_hd__or2_1 _3369_ (.A(net297),
    .B(_0744_),
    .X(_0813_));
 sky130_fd_sc_hd__nand2_1 _3370_ (.A(_0745_),
    .B(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__a311o_1 _3371_ (.A1(_0749_),
    .A2(_0752_),
    .A3(_0811_),
    .B1(_0812_),
    .C1(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__nor2_1 _3372_ (.A(net295),
    .B(_0741_),
    .Y(_0816_));
 sky130_fd_sc_hd__or2_1 _3373_ (.A(_0742_),
    .B(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__a21oi_2 _3374_ (.A1(_0745_),
    .A2(_0815_),
    .B1(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__nor2_1 _3375_ (.A(net293),
    .B(_0729_),
    .Y(_0819_));
 sky130_fd_sc_hd__or2_1 _3376_ (.A(_0730_),
    .B(_0819_),
    .X(_0820_));
 sky130_fd_sc_hd__or2_1 _3377_ (.A(_0726_),
    .B(_0727_),
    .X(_0821_));
 sky130_fd_sc_hd__nor3_1 _3378_ (.A(_0723_),
    .B(_0820_),
    .C(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__o211ai_2 _3379_ (.A1(_0742_),
    .A2(_0818_),
    .B1(_0822_),
    .C1(_0714_),
    .Y(_0823_));
 sky130_fd_sc_hd__xor2_2 _3380_ (.A(_0654_),
    .B(_0660_),
    .X(_0824_));
 sky130_fd_sc_hd__xnor2_1 _3381_ (.A(net269),
    .B(_0824_),
    .Y(_0825_));
 sky130_fd_sc_hd__o21ai_1 _3382_ (.A1(_0481_),
    .A2(_0649_),
    .B1(_1928_),
    .Y(_0826_));
 sky130_fd_sc_hd__xnor2_2 _3383_ (.A(_0653_),
    .B(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__xnor2_2 _3384_ (.A(net271),
    .B(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__a31o_1 _3385_ (.A1(_0631_),
    .A2(_0636_),
    .A3(_0643_),
    .B1(_0701_),
    .X(_0829_));
 sky130_fd_sc_hd__xor2_1 _3386_ (.A(_0648_),
    .B(_0829_),
    .X(_0830_));
 sky130_fd_sc_hd__nand2_1 _3387_ (.A(net276),
    .B(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__or2_1 _3388_ (.A(net276),
    .B(_0830_),
    .X(_0832_));
 sky130_fd_sc_hd__nand2_1 _3389_ (.A(_0831_),
    .B(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__a21o_1 _3390_ (.A1(_0648_),
    .A2(_0829_),
    .B1(_0668_),
    .X(_0834_));
 sky130_fd_sc_hd__xnor2_2 _3391_ (.A(_0481_),
    .B(_0834_),
    .Y(_0835_));
 sky130_fd_sc_hd__xor2_1 _3392_ (.A(net273),
    .B(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__or4b_1 _3393_ (.A(_0825_),
    .B(_0828_),
    .C(_0833_),
    .D_N(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__a21oi_1 _3394_ (.A1(_0737_),
    .A2(_0823_),
    .B1(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__nand2_1 _3395_ (.A(net273),
    .B(_0835_),
    .Y(_0839_));
 sky130_fd_sc_hd__nor2_1 _3396_ (.A(net273),
    .B(_0835_),
    .Y(_0840_));
 sky130_fd_sc_hd__a2111oi_1 _3397_ (.A1(_0831_),
    .A2(_0839_),
    .B1(_0840_),
    .C1(_0825_),
    .D1(_0828_),
    .Y(_0841_));
 sky130_fd_sc_hd__a22o_1 _3398_ (.A1(net269),
    .A2(_0824_),
    .B1(_0827_),
    .B2(net271),
    .X(_0842_));
 sky130_fd_sc_hd__o21a_1 _3399_ (.A1(net270),
    .A2(_0824_),
    .B1(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__xnor2_1 _3400_ (.A(net268),
    .B(_0692_),
    .Y(_0844_));
 sky130_fd_sc_hd__o31ai_2 _3401_ (.A1(_0838_),
    .A2(net260),
    .A3(_0843_),
    .B1(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__xnor2_1 _3402_ (.A(_0670_),
    .B(_0471_),
    .Y(_0846_));
 sky130_fd_sc_hd__nand2_1 _3403_ (.A(net267),
    .B(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__nor2_1 _3404_ (.A(net267),
    .B(_0846_),
    .Y(_0848_));
 sky130_fd_sc_hd__a31o_1 _3405_ (.A1(_0693_),
    .A2(_0845_),
    .A3(_0847_),
    .B1(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__or2_1 _3406_ (.A(_0690_),
    .B(_0849_),
    .X(_0850_));
 sky130_fd_sc_hd__o31a_2 _3407_ (.A1(_2158_),
    .A2(_0682_),
    .A3(_0683_),
    .B1(_0680_),
    .X(_0851_));
 sky130_fd_sc_hd__a221o_1 _3408_ (.A1(_1942_),
    .A2(net187),
    .B1(_1966_),
    .B2(net117),
    .C1(_1952_),
    .X(_0852_));
 sky130_fd_sc_hd__a21o_1 _3409_ (.A1(net152),
    .A2(_1946_),
    .B1(_0852_),
    .X(_0853_));
 sky130_fd_sc_hd__o21ai_2 _3410_ (.A1(net95),
    .A2(_1935_),
    .B1(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__xnor2_4 _3411_ (.A(\sum[31] ),
    .B(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__xnor2_4 _3412_ (.A(_0851_),
    .B(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__a21bo_1 _3413_ (.A1(_0673_),
    .A2(_0675_),
    .B1_N(_0672_),
    .X(_0857_));
 sky130_fd_sc_hd__xnor2_2 _3414_ (.A(\workunit2[31] ),
    .B(\workunit1[31] ),
    .Y(_0858_));
 sky130_fd_sc_hd__xor2_1 _3415_ (.A(net327),
    .B(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__xnor2_1 _3416_ (.A(_0857_),
    .B(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__xnor2_1 _3417_ (.A(_0856_),
    .B(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__o21ba_1 _3418_ (.A1(_0669_),
    .A2(_0686_),
    .B1_N(_0671_),
    .X(_0862_));
 sky130_fd_sc_hd__xnor2_1 _3419_ (.A(_0861_),
    .B(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__a21o_1 _3420_ (.A1(_0688_),
    .A2(_0850_),
    .B1(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__nand3_1 _3421_ (.A(_0688_),
    .B(_0850_),
    .C(_0863_),
    .Y(_0865_));
 sky130_fd_sc_hd__inv_2 _3422_ (.A(net262),
    .Y(_0866_));
 sky130_fd_sc_hd__buf_1 _3423_ (.A(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__inv_2 _3424_ (.A(\state[0] ),
    .Y(_0868_));
 sky130_fd_sc_hd__or2_1 _3425_ (.A(\state[4] ),
    .B(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3426_ (.A(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__nor2_1 _3427_ (.A(net264),
    .B(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__and3_2 _3428_ (.A(_0867_),
    .B(_0769_),
    .C(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3429_ (.A(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__buf_4 _3430_ (.A(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__nor2_1 _3431_ (.A(_1923_),
    .B(_0872_),
    .Y(_0875_));
 sky130_fd_sc_hd__buf_2 _3432_ (.A(_0875_),
    .X(_0876_));
 sky130_fd_sc_hd__a22o_1 _3433_ (.A1(net483),
    .A2(_0874_),
    .B1(_0876_),
    .B2(\workunit2[31] ),
    .X(_0877_));
 sky130_fd_sc_hd__a31o_1 _3434_ (.A1(_1926_),
    .A2(_0864_),
    .A3(_0865_),
    .B1(_0877_),
    .X(_0352_));
 sky130_fd_sc_hd__buf_2 _3435_ (.A(_1924_),
    .X(_0878_));
 sky130_fd_sc_hd__nand2_1 _3436_ (.A(_0690_),
    .B(_0849_),
    .Y(_0879_));
 sky130_fd_sc_hd__clkbuf_4 _3437_ (.A(_0873_),
    .X(_0880_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3438_ (.A(_0875_),
    .X(_0881_));
 sky130_fd_sc_hd__buf_2 _3439_ (.A(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__a22o_1 _3440_ (.A1(net490),
    .A2(_0880_),
    .B1(_0882_),
    .B2(\workunit2[30] ),
    .X(_0883_));
 sky130_fd_sc_hd__a31o_1 _3441_ (.A1(_0878_),
    .A2(_0850_),
    .A3(_0879_),
    .B1(_0883_),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_2 _3442_ (.A(_0881_),
    .X(_0884_));
 sky130_fd_sc_hd__and2b_1 _3443_ (.A_N(_0848_),
    .B(_0847_),
    .X(_0885_));
 sky130_fd_sc_hd__a21oi_1 _3444_ (.A1(_0693_),
    .A2(_0845_),
    .B1(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__a31o_1 _3445_ (.A1(_0693_),
    .A2(_0845_),
    .A3(_0885_),
    .B1(_0513_),
    .X(_0887_));
 sky130_fd_sc_hd__or2_1 _3446_ (.A(_0886_),
    .B(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__clkbuf_4 _3447_ (.A(_0873_),
    .X(_0889_));
 sky130_fd_sc_hd__a21o_1 _3448_ (.A1(net510),
    .A2(_0889_),
    .B1(_1925_),
    .X(_0890_));
 sky130_fd_sc_hd__a22o_1 _3449_ (.A1(\workunit2[29] ),
    .A2(_0884_),
    .B1(_0888_),
    .B2(_0890_),
    .X(_0350_));
 sky130_fd_sc_hd__or4_1 _3450_ (.A(_0844_),
    .B(_0838_),
    .C(_0841_),
    .D(_0843_),
    .X(_0891_));
 sky130_fd_sc_hd__a22o_1 _3451_ (.A1(net522),
    .A2(_0880_),
    .B1(_0876_),
    .B2(net268),
    .X(_0892_));
 sky130_fd_sc_hd__a31o_1 _3452_ (.A1(_1926_),
    .A2(_0845_),
    .A3(_0891_),
    .B1(_0892_),
    .X(_0349_));
 sky130_fd_sc_hd__buf_2 _3453_ (.A(_0872_),
    .X(_0893_));
 sky130_fd_sc_hd__buf_2 _3454_ (.A(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__clkbuf_2 _3455_ (.A(_0881_),
    .X(_0895_));
 sky130_fd_sc_hd__clkbuf_2 _3456_ (.A(_0513_),
    .X(_0896_));
 sky130_fd_sc_hd__a21o_1 _3457_ (.A1(_0737_),
    .A2(_0823_),
    .B1(_0833_),
    .X(_0897_));
 sky130_fd_sc_hd__a31o_1 _3458_ (.A1(_0831_),
    .A2(_0839_),
    .A3(_0897_),
    .B1(_0840_),
    .X(_0898_));
 sky130_fd_sc_hd__o2bb2a_1 _3459_ (.A1_N(net271),
    .A2_N(_0827_),
    .B1(_0828_),
    .B2(_0898_),
    .X(_0899_));
 sky130_fd_sc_hd__xnor2_1 _3460_ (.A(_0825_),
    .B(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__nor2_1 _3461_ (.A(_0896_),
    .B(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__a221o_1 _3462_ (.A1(net473),
    .A2(_0894_),
    .B1(_0895_),
    .B2(net269),
    .C1(_0901_),
    .X(_0348_));
 sky130_fd_sc_hd__buf_2 _3463_ (.A(_0893_),
    .X(_0902_));
 sky130_fd_sc_hd__o21a_1 _3464_ (.A1(_0828_),
    .A2(_0898_),
    .B1(_1924_),
    .X(_0903_));
 sky130_fd_sc_hd__a21boi_1 _3465_ (.A1(_0828_),
    .A2(_0898_),
    .B1_N(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__a221o_1 _3466_ (.A1(net465),
    .A2(_0902_),
    .B1(_0895_),
    .B2(net271),
    .C1(_0904_),
    .X(_0347_));
 sky130_fd_sc_hd__nand2_1 _3467_ (.A(_0831_),
    .B(_0897_),
    .Y(_0905_));
 sky130_fd_sc_hd__xor2_1 _3468_ (.A(_0836_),
    .B(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__clkbuf_2 _3469_ (.A(_0873_),
    .X(_0907_));
 sky130_fd_sc_hd__clkbuf_2 _3470_ (.A(_0881_),
    .X(_0908_));
 sky130_fd_sc_hd__a22o_1 _3471_ (.A1(net492),
    .A2(_0907_),
    .B1(_0908_),
    .B2(net275),
    .X(_0909_));
 sky130_fd_sc_hd__a21o_1 _3472_ (.A1(_0878_),
    .A2(_0906_),
    .B1(_0909_),
    .X(_0346_));
 sky130_fd_sc_hd__buf_2 _3473_ (.A(_1924_),
    .X(_0910_));
 sky130_fd_sc_hd__nand3_1 _3474_ (.A(_0737_),
    .B(_0823_),
    .C(_0833_),
    .Y(_0911_));
 sky130_fd_sc_hd__a22o_1 _3475_ (.A1(net551),
    .A2(_0880_),
    .B1(_0882_),
    .B2(net277),
    .X(_0912_));
 sky130_fd_sc_hd__a31o_1 _3476_ (.A1(_0910_),
    .A2(_0897_),
    .A3(_0911_),
    .B1(_0912_),
    .X(_0345_));
 sky130_fd_sc_hd__inv_2 _3477_ (.A(_0734_),
    .Y(_0913_));
 sky130_fd_sc_hd__o21ai_1 _3478_ (.A1(_0742_),
    .A2(_0818_),
    .B1(_0822_),
    .Y(_0914_));
 sky130_fd_sc_hd__a21boi_1 _3479_ (.A1(_0913_),
    .A2(_0914_),
    .B1_N(_0712_),
    .Y(_0915_));
 sky130_fd_sc_hd__nor3_1 _3480_ (.A(_0704_),
    .B(_0708_),
    .C(_0915_),
    .Y(_0916_));
 sky130_fd_sc_hd__nand2_1 _3481_ (.A(net280),
    .B(_0698_),
    .Y(_0917_));
 sky130_fd_sc_hd__o31a_1 _3482_ (.A1(_0699_),
    .A2(_0709_),
    .A3(_0916_),
    .B1(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__xnor2_1 _3483_ (.A(_0696_),
    .B(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__nand2_1 _3484_ (.A(_0910_),
    .B(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__a21o_1 _3485_ (.A1(net500),
    .A2(_0889_),
    .B1(_1925_),
    .X(_0921_));
 sky130_fd_sc_hd__a22o_1 _3486_ (.A1(net279),
    .A2(_0884_),
    .B1(_0920_),
    .B2(_0921_),
    .X(_0344_));
 sky130_fd_sc_hd__o21ai_1 _3487_ (.A1(_0709_),
    .A2(_0916_),
    .B1(_0699_),
    .Y(_0922_));
 sky130_fd_sc_hd__o31a_1 _3488_ (.A1(_0699_),
    .A2(_0709_),
    .A3(_0916_),
    .B1(_0910_),
    .X(_0923_));
 sky130_fd_sc_hd__a22o_1 _3489_ (.A1(net486),
    .A2(_0907_),
    .B1(_0908_),
    .B2(net280),
    .X(_0924_));
 sky130_fd_sc_hd__a21o_1 _3490_ (.A1(_0922_),
    .A2(_0923_),
    .B1(_0924_),
    .X(_0343_));
 sky130_fd_sc_hd__nor2_1 _3491_ (.A(_0704_),
    .B(_0915_),
    .Y(_0925_));
 sky130_fd_sc_hd__xnor2_1 _3492_ (.A(_0713_),
    .B(_0925_),
    .Y(_0926_));
 sky130_fd_sc_hd__mux2_1 _3493_ (.A0(net565),
    .A1(_0926_),
    .S(_1923_),
    .X(_0927_));
 sky130_fd_sc_hd__mux2_1 _3494_ (.A0(_0927_),
    .A1(net282),
    .S(_0881_),
    .X(_0928_));
 sky130_fd_sc_hd__clkbuf_1 _3495_ (.A(_0928_),
    .X(_0342_));
 sky130_fd_sc_hd__or3b_1 _3496_ (.A(_0712_),
    .B(_0734_),
    .C_N(_0914_),
    .X(_0929_));
 sky130_fd_sc_hd__nor2_1 _3497_ (.A(_0896_),
    .B(_0915_),
    .Y(_0930_));
 sky130_fd_sc_hd__a22o_1 _3498_ (.A1(net481),
    .A2(_0907_),
    .B1(_0908_),
    .B2(net284),
    .X(_0931_));
 sky130_fd_sc_hd__a21o_1 _3499_ (.A1(_0929_),
    .A2(_0930_),
    .B1(_0931_),
    .X(_0341_));
 sky130_fd_sc_hd__a21o_1 _3500_ (.A1(net496),
    .A2(_0907_),
    .B1(_1925_),
    .X(_0932_));
 sky130_fd_sc_hd__o21bai_1 _3501_ (.A1(_0742_),
    .A2(_0818_),
    .B1_N(_0820_),
    .Y(_0933_));
 sky130_fd_sc_hd__and2_1 _3502_ (.A(_0731_),
    .B(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__or3_1 _3503_ (.A(_0722_),
    .B(_0726_),
    .C(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__a21oi_1 _3504_ (.A1(_0720_),
    .A2(_0935_),
    .B1(_0717_),
    .Y(_0936_));
 sky130_fd_sc_hd__and3_1 _3505_ (.A(_0717_),
    .B(_0720_),
    .C(_0935_),
    .X(_0937_));
 sky130_fd_sc_hd__o21ai_1 _3506_ (.A1(_0936_),
    .A2(_0937_),
    .B1(_0910_),
    .Y(_0938_));
 sky130_fd_sc_hd__a22o_1 _3507_ (.A1(net288),
    .A2(_0884_),
    .B1(_0932_),
    .B2(_0938_),
    .X(_0340_));
 sky130_fd_sc_hd__o21ai_1 _3508_ (.A1(_0726_),
    .A2(_0934_),
    .B1(_0722_),
    .Y(_0939_));
 sky130_fd_sc_hd__clkbuf_2 _3509_ (.A(_0873_),
    .X(_0940_));
 sky130_fd_sc_hd__a22o_1 _3510_ (.A1(net513),
    .A2(_0940_),
    .B1(_0882_),
    .B2(net290),
    .X(_0941_));
 sky130_fd_sc_hd__a31o_1 _3511_ (.A1(_0910_),
    .A2(_0935_),
    .A3(_0939_),
    .B1(_0941_),
    .X(_0339_));
 sky130_fd_sc_hd__or2b_1 _3512_ (.A(_0730_),
    .B_N(_0933_),
    .X(_0942_));
 sky130_fd_sc_hd__xnor2_1 _3513_ (.A(_0821_),
    .B(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__mux2_1 _3514_ (.A0(net573),
    .A1(_0943_),
    .S(_1923_),
    .X(_0944_));
 sky130_fd_sc_hd__mux2_1 _3515_ (.A0(_0944_),
    .A1(net292),
    .S(_0876_),
    .X(_0945_));
 sky130_fd_sc_hd__clkbuf_1 _3516_ (.A(_0945_),
    .X(_0338_));
 sky130_fd_sc_hd__or3b_1 _3517_ (.A(_0742_),
    .B(_0818_),
    .C_N(_0820_),
    .X(_0946_));
 sky130_fd_sc_hd__a22o_1 _3518_ (.A1(net508),
    .A2(_0874_),
    .B1(_0882_),
    .B2(net294),
    .X(_0947_));
 sky130_fd_sc_hd__a31o_1 _3519_ (.A1(_0878_),
    .A2(_0933_),
    .A3(_0946_),
    .B1(_0947_),
    .X(_0337_));
 sky130_fd_sc_hd__and3_1 _3520_ (.A(_0817_),
    .B(_0745_),
    .C(_0815_),
    .X(_0948_));
 sky130_fd_sc_hd__buf_2 _3521_ (.A(_0893_),
    .X(_0949_));
 sky130_fd_sc_hd__a22oi_1 _3522_ (.A1(net471),
    .A2(_0949_),
    .B1(_0895_),
    .B2(net296),
    .Y(_0950_));
 sky130_fd_sc_hd__o31ai_1 _3523_ (.A1(_0896_),
    .A2(_0818_),
    .A3(_0948_),
    .B1(_0950_),
    .Y(_0336_));
 sky130_fd_sc_hd__a31o_1 _3524_ (.A1(_0749_),
    .A2(_0752_),
    .A3(_0811_),
    .B1(_0812_),
    .X(_0951_));
 sky130_fd_sc_hd__nand2_1 _3525_ (.A(_1924_),
    .B(_0815_),
    .Y(_0952_));
 sky130_fd_sc_hd__a21oi_1 _3526_ (.A1(_0814_),
    .A2(_0951_),
    .B1(_0952_),
    .Y(_0953_));
 sky130_fd_sc_hd__a221o_1 _3527_ (.A1(net469),
    .A2(_0902_),
    .B1(_0895_),
    .B2(net298),
    .C1(_0953_),
    .X(_0335_));
 sky130_fd_sc_hd__and2_1 _3528_ (.A(_0752_),
    .B(_0811_),
    .X(_0954_));
 sky130_fd_sc_hd__and2b_1 _3529_ (.A_N(_0812_),
    .B(_0749_),
    .X(_0955_));
 sky130_fd_sc_hd__a21oi_1 _3530_ (.A1(_0954_),
    .A2(_0955_),
    .B1(_0513_),
    .Y(_0956_));
 sky130_fd_sc_hd__o21ai_1 _3531_ (.A1(_0954_),
    .A2(_0955_),
    .B1(_0956_),
    .Y(_0957_));
 sky130_fd_sc_hd__a21o_1 _3532_ (.A1(net520),
    .A2(_0889_),
    .B1(_1925_),
    .X(_0958_));
 sky130_fd_sc_hd__a22o_1 _3533_ (.A1(net300),
    .A2(_0884_),
    .B1(_0957_),
    .B2(_0958_),
    .X(_0334_));
 sky130_fd_sc_hd__a31o_1 _3534_ (.A1(_0755_),
    .A2(_0757_),
    .A3(_0808_),
    .B1(_0809_),
    .X(_0959_));
 sky130_fd_sc_hd__nand2_1 _3535_ (.A(_0810_),
    .B(_0959_),
    .Y(_0960_));
 sky130_fd_sc_hd__and3_1 _3536_ (.A(_1924_),
    .B(_0811_),
    .C(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__a22o_1 _3537_ (.A1(net582),
    .A2(_0873_),
    .B1(_0881_),
    .B2(net302),
    .X(_0962_));
 sky130_fd_sc_hd__or2_1 _3538_ (.A(_0961_),
    .B(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__clkbuf_1 _3539_ (.A(_0963_),
    .X(_0333_));
 sky130_fd_sc_hd__and2_1 _3540_ (.A(_0757_),
    .B(_0808_),
    .X(_0964_));
 sky130_fd_sc_hd__or2b_1 _3541_ (.A(_0809_),
    .B_N(_0755_),
    .X(_0965_));
 sky130_fd_sc_hd__xnor2_1 _3542_ (.A(_0964_),
    .B(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__nor2_1 _3543_ (.A(_0896_),
    .B(_0966_),
    .Y(_0967_));
 sky130_fd_sc_hd__a221o_1 _3544_ (.A1(net463),
    .A2(_0902_),
    .B1(_0884_),
    .B2(net304),
    .C1(_0967_),
    .X(_0332_));
 sky130_fd_sc_hd__a31o_1 _3545_ (.A1(_0760_),
    .A2(_0762_),
    .A3(_0803_),
    .B1(_0804_),
    .X(_0968_));
 sky130_fd_sc_hd__nand2_1 _3546_ (.A(_0807_),
    .B(_0968_),
    .Y(_0969_));
 sky130_fd_sc_hd__and2_1 _3547_ (.A(_0808_),
    .B(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__a22o_1 _3548_ (.A1(net575),
    .A2(_0889_),
    .B1(_0908_),
    .B2(net306),
    .X(_0971_));
 sky130_fd_sc_hd__a21o_1 _3549_ (.A1(_0878_),
    .A2(_0970_),
    .B1(_0971_),
    .X(_0331_));
 sky130_fd_sc_hd__a21o_1 _3550_ (.A1(net502),
    .A2(_0907_),
    .B1(_1925_),
    .X(_0972_));
 sky130_fd_sc_hd__or2_1 _3551_ (.A(net307),
    .B(_0759_),
    .X(_0973_));
 sky130_fd_sc_hd__and4_1 _3552_ (.A(_0760_),
    .B(_0973_),
    .C(_0762_),
    .D(_0803_),
    .X(_0974_));
 sky130_fd_sc_hd__a22o_1 _3553_ (.A1(_0760_),
    .A2(_0973_),
    .B1(_0762_),
    .B2(_0803_),
    .X(_0975_));
 sky130_fd_sc_hd__or3b_1 _3554_ (.A(_0513_),
    .B(_0974_),
    .C_N(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__a22o_1 _3555_ (.A1(net308),
    .A2(_0884_),
    .B1(_0972_),
    .B2(_0976_),
    .X(_0330_));
 sky130_fd_sc_hd__or3_1 _3556_ (.A(_0765_),
    .B(_0800_),
    .C(_0802_),
    .X(_0977_));
 sky130_fd_sc_hd__a22o_1 _3557_ (.A1(net571),
    .A2(_0880_),
    .B1(_0882_),
    .B2(net309),
    .X(_0978_));
 sky130_fd_sc_hd__a31o_1 _3558_ (.A1(_1926_),
    .A2(_0803_),
    .A3(_0977_),
    .B1(_0978_),
    .X(_0329_));
 sky130_fd_sc_hd__and3_1 _3559_ (.A(_0799_),
    .B(_0768_),
    .C(_0797_),
    .X(_0979_));
 sky130_fd_sc_hd__a22oi_1 _3560_ (.A1(net526),
    .A2(_0949_),
    .B1(_0895_),
    .B2(net311),
    .Y(_0980_));
 sky130_fd_sc_hd__o31ai_1 _3561_ (.A1(_0896_),
    .A2(_0800_),
    .A3(_0979_),
    .B1(_0980_),
    .Y(_0328_));
 sky130_fd_sc_hd__nor2_1 _3562_ (.A(_0772_),
    .B(_0795_),
    .Y(_0981_));
 sky130_fd_sc_hd__nand2_1 _3563_ (.A(_0796_),
    .B(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__a22o_1 _3564_ (.A1(net535),
    .A2(_0940_),
    .B1(_0908_),
    .B2(net314),
    .X(_0983_));
 sky130_fd_sc_hd__a31o_1 _3565_ (.A1(_1926_),
    .A2(_0797_),
    .A3(_0982_),
    .B1(_0983_),
    .X(_0327_));
 sky130_fd_sc_hd__and3_1 _3566_ (.A(_0794_),
    .B(_0774_),
    .C(_0793_),
    .X(_0984_));
 sky130_fd_sc_hd__nor3_1 _3567_ (.A(_0896_),
    .B(_0795_),
    .C(_0984_),
    .Y(_0985_));
 sky130_fd_sc_hd__a221o_1 _3568_ (.A1(net506),
    .A2(_0902_),
    .B1(_0895_),
    .B2(net316),
    .C1(_0985_),
    .X(_0326_));
 sky130_fd_sc_hd__nand3_1 _3569_ (.A(_0776_),
    .B(_0791_),
    .C(_0792_),
    .Y(_0986_));
 sky130_fd_sc_hd__a22o_1 _3570_ (.A1(net524),
    .A2(_0940_),
    .B1(_0876_),
    .B2(\workunit2[4] ),
    .X(_0987_));
 sky130_fd_sc_hd__a31o_1 _3571_ (.A1(_1926_),
    .A2(_0793_),
    .A3(_0986_),
    .B1(_0987_),
    .X(_0325_));
 sky130_fd_sc_hd__nand3_1 _3572_ (.A(_0790_),
    .B(_0779_),
    .C(_0789_),
    .Y(_0988_));
 sky130_fd_sc_hd__a22o_1 _3573_ (.A1(net580),
    .A2(_0940_),
    .B1(_0876_),
    .B2(\workunit2[3] ),
    .X(_0989_));
 sky130_fd_sc_hd__a31o_1 _3574_ (.A1(_1926_),
    .A2(_0791_),
    .A3(_0988_),
    .B1(_0989_),
    .X(_0324_));
 sky130_fd_sc_hd__o21ai_1 _3575_ (.A1(_0780_),
    .A2(_0788_),
    .B1(_0787_),
    .Y(_0990_));
 sky130_fd_sc_hd__a22o_1 _3576_ (.A1(net584),
    .A2(_0940_),
    .B1(_0882_),
    .B2(net320),
    .X(_0991_));
 sky130_fd_sc_hd__a31o_1 _3577_ (.A1(_0878_),
    .A2(_0789_),
    .A3(_0990_),
    .B1(_0991_),
    .X(_0323_));
 sky130_fd_sc_hd__nor2_1 _3578_ (.A(_0786_),
    .B(_0785_),
    .Y(_0992_));
 sky130_fd_sc_hd__xnor2_1 _3579_ (.A(_0781_),
    .B(_0992_),
    .Y(_0993_));
 sky130_fd_sc_hd__a22o_1 _3580_ (.A1(net528),
    .A2(_0907_),
    .B1(_0908_),
    .B2(\workunit2[1] ),
    .X(_0994_));
 sky130_fd_sc_hd__a21o_1 _3581_ (.A1(_0878_),
    .A2(_0993_),
    .B1(_0994_),
    .X(_0322_));
 sky130_fd_sc_hd__or2_1 _3582_ (.A(\workunit2[0] ),
    .B(_0554_),
    .X(_0995_));
 sky130_fd_sc_hd__a22o_1 _3583_ (.A1(net577),
    .A2(_0940_),
    .B1(_0876_),
    .B2(net322),
    .X(_0996_));
 sky130_fd_sc_hd__a31o_1 _3584_ (.A1(_0910_),
    .A2(_0781_),
    .A3(_0995_),
    .B1(_0996_),
    .X(_0321_));
 sky130_fd_sc_hd__inv_2 _3585_ (.A(net264),
    .Y(_0997_));
 sky130_fd_sc_hd__nand2_1 _3586_ (.A(_0866_),
    .B(net261),
    .Y(_0998_));
 sky130_fd_sc_hd__or2_2 _3587_ (.A(_0870_),
    .B(_0998_),
    .X(_0999_));
 sky130_fd_sc_hd__nor2_1 _3588_ (.A(_0997_),
    .B(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__buf_1 _3589_ (.A(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__buf_2 _3590_ (.A(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__nand2_1 _3591_ (.A(net269),
    .B(net278),
    .Y(_1003_));
 sky130_fd_sc_hd__or2_1 _3592_ (.A(net270),
    .B(net278),
    .X(_1004_));
 sky130_fd_sc_hd__nand2_1 _3593_ (.A(_1003_),
    .B(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__xor2_1 _3594_ (.A(\workunit2[31] ),
    .B(net281),
    .X(_1006_));
 sky130_fd_sc_hd__nand2_1 _3595_ (.A(net272),
    .B(_1006_),
    .Y(_1007_));
 sky130_fd_sc_hd__or2_1 _3596_ (.A(net266),
    .B(net283),
    .X(_1008_));
 sky130_fd_sc_hd__nand2_1 _3597_ (.A(net266),
    .B(net283),
    .Y(_1009_));
 sky130_fd_sc_hd__nand3_1 _3598_ (.A(net273),
    .B(_1008_),
    .C(_1009_),
    .Y(_1010_));
 sky130_fd_sc_hd__or2_1 _3599_ (.A(net267),
    .B(net285),
    .X(_1011_));
 sky130_fd_sc_hd__nand2_1 _3600_ (.A(net267),
    .B(net285),
    .Y(_1012_));
 sky130_fd_sc_hd__a21o_1 _3601_ (.A1(_1011_),
    .A2(_1012_),
    .B1(net276),
    .X(_1013_));
 sky130_fd_sc_hd__or2_1 _3602_ (.A(net268),
    .B(net286),
    .X(_1014_));
 sky130_fd_sc_hd__nand2_1 _3603_ (.A(net268),
    .B(net287),
    .Y(_1015_));
 sky130_fd_sc_hd__nand3_1 _3604_ (.A(net278),
    .B(_1014_),
    .C(_1015_),
    .Y(_1016_));
 sky130_fd_sc_hd__or2_1 _3605_ (.A(net269),
    .B(net289),
    .X(_1017_));
 sky130_fd_sc_hd__nand2_1 _3606_ (.A(net269),
    .B(net290),
    .Y(_1018_));
 sky130_fd_sc_hd__nand3_1 _3607_ (.A(net280),
    .B(_1017_),
    .C(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__a21oi_1 _3608_ (.A1(_1014_),
    .A2(_1015_),
    .B1(net278),
    .Y(_1020_));
 sky130_fd_sc_hd__a21oi_1 _3609_ (.A1(_1016_),
    .A2(_1019_),
    .B1(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__xor2_1 _3610_ (.A(net275),
    .B(net293),
    .X(_1022_));
 sky130_fd_sc_hd__nand2_1 _3611_ (.A(net284),
    .B(_1022_),
    .Y(_1023_));
 sky130_fd_sc_hd__or2_1 _3612_ (.A(net271),
    .B(net291),
    .X(_1024_));
 sky130_fd_sc_hd__nand2_1 _3613_ (.A(net271),
    .B(net291),
    .Y(_1025_));
 sky130_fd_sc_hd__nand3_1 _3614_ (.A(net282),
    .B(_1024_),
    .C(_1025_),
    .Y(_1026_));
 sky130_fd_sc_hd__a21oi_1 _3615_ (.A1(_1024_),
    .A2(_1025_),
    .B1(net282),
    .Y(_1027_));
 sky130_fd_sc_hd__a21oi_1 _3616_ (.A1(_1023_),
    .A2(_1026_),
    .B1(_1027_),
    .Y(_1028_));
 sky130_fd_sc_hd__or2_1 _3617_ (.A(net277),
    .B(net295),
    .X(_1029_));
 sky130_fd_sc_hd__nand2_1 _3618_ (.A(net277),
    .B(net295),
    .Y(_1030_));
 sky130_fd_sc_hd__a21oi_1 _3619_ (.A1(_1029_),
    .A2(_1030_),
    .B1(net286),
    .Y(_1031_));
 sky130_fd_sc_hd__inv_2 _3620_ (.A(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__or2_1 _3621_ (.A(net278),
    .B(net297),
    .X(_1033_));
 sky130_fd_sc_hd__nand2_1 _3622_ (.A(net278),
    .B(net297),
    .Y(_1034_));
 sky130_fd_sc_hd__and3_1 _3623_ (.A(net289),
    .B(_1033_),
    .C(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__a32o_1 _3624_ (.A1(net286),
    .A2(_1029_),
    .A3(_1030_),
    .B1(_1032_),
    .B2(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__or2_1 _3625_ (.A(net284),
    .B(net303),
    .X(_1037_));
 sky130_fd_sc_hd__nand2_1 _3626_ (.A(net284),
    .B(net303),
    .Y(_1038_));
 sky130_fd_sc_hd__a21o_1 _3627_ (.A1(_1037_),
    .A2(_1038_),
    .B1(net295),
    .X(_1039_));
 sky130_fd_sc_hd__or2_1 _3628_ (.A(net286),
    .B(net306),
    .X(_1040_));
 sky130_fd_sc_hd__nand2_1 _3629_ (.A(net286),
    .B(net305),
    .Y(_1041_));
 sky130_fd_sc_hd__a21o_1 _3630_ (.A1(_1040_),
    .A2(_1041_),
    .B1(net298),
    .X(_1042_));
 sky130_fd_sc_hd__nand3_1 _3631_ (.A(net295),
    .B(_1037_),
    .C(_1038_),
    .Y(_1043_));
 sky130_fd_sc_hd__a21boi_1 _3632_ (.A1(_1039_),
    .A2(_1042_),
    .B1_N(_1043_),
    .Y(_1044_));
 sky130_fd_sc_hd__inv_2 _3633_ (.A(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__or2_1 _3634_ (.A(net301),
    .B(net318),
    .X(_1046_));
 sky130_fd_sc_hd__nand2_1 _3635_ (.A(net301),
    .B(net318),
    .Y(_1047_));
 sky130_fd_sc_hd__a21o_1 _3636_ (.A1(_1046_),
    .A2(_1047_),
    .B1(net311),
    .X(_1048_));
 sky130_fd_sc_hd__or2_1 _3637_ (.A(net303),
    .B(net319),
    .X(_1049_));
 sky130_fd_sc_hd__nand2_1 _3638_ (.A(net303),
    .B(net320),
    .Y(_1050_));
 sky130_fd_sc_hd__a21o_1 _3639_ (.A1(_1049_),
    .A2(_1050_),
    .B1(net313),
    .X(_1051_));
 sky130_fd_sc_hd__or2_1 _3640_ (.A(net309),
    .B(net318),
    .X(_1052_));
 sky130_fd_sc_hd__xor2_2 _3641_ (.A(net313),
    .B(net321),
    .X(_1053_));
 sky130_fd_sc_hd__and2_1 _3642_ (.A(net313),
    .B(net321),
    .X(_1054_));
 sky130_fd_sc_hd__a31o_1 _3643_ (.A1(net315),
    .A2(net322),
    .A3(_1053_),
    .B1(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__or2_1 _3644_ (.A(net311),
    .B(net319),
    .X(_1056_));
 sky130_fd_sc_hd__nand2_1 _3645_ (.A(net311),
    .B(net319),
    .Y(_1057_));
 sky130_fd_sc_hd__a21bo_1 _3646_ (.A1(_1055_),
    .A2(_1056_),
    .B1_N(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__nand2_1 _3647_ (.A(net309),
    .B(net318),
    .Y(_1059_));
 sky130_fd_sc_hd__a21bo_1 _3648_ (.A1(_1052_),
    .A2(_1058_),
    .B1_N(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__xor2_1 _3649_ (.A(net307),
    .B(net322),
    .X(_1061_));
 sky130_fd_sc_hd__xnor2_1 _3650_ (.A(net317),
    .B(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__or2_1 _3651_ (.A(net305),
    .B(net321),
    .X(_1063_));
 sky130_fd_sc_hd__nand2_1 _3652_ (.A(net305),
    .B(net321),
    .Y(_1064_));
 sky130_fd_sc_hd__a21oi_1 _3653_ (.A1(_1063_),
    .A2(_1064_),
    .B1(net315),
    .Y(_1065_));
 sky130_fd_sc_hd__and3_1 _3654_ (.A(net315),
    .B(_1063_),
    .C(_1064_),
    .X(_1066_));
 sky130_fd_sc_hd__or2_1 _3655_ (.A(_1065_),
    .B(_1066_),
    .X(_1067_));
 sky130_fd_sc_hd__nor2_1 _3656_ (.A(_1062_),
    .B(_1067_),
    .Y(_1068_));
 sky130_fd_sc_hd__and3b_1 _3657_ (.A_N(_1065_),
    .B(_1061_),
    .C(net317),
    .X(_1069_));
 sky130_fd_sc_hd__a211o_1 _3658_ (.A1(_1060_),
    .A2(_1068_),
    .B1(_1069_),
    .C1(_1066_),
    .X(_1070_));
 sky130_fd_sc_hd__and3_1 _3659_ (.A(net313),
    .B(_1049_),
    .C(_1050_),
    .X(_1071_));
 sky130_fd_sc_hd__a21o_1 _3660_ (.A1(_1051_),
    .A2(_1070_),
    .B1(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__and3_1 _3661_ (.A(net311),
    .B(_1046_),
    .C(_1047_),
    .X(_1073_));
 sky130_fd_sc_hd__a21o_1 _3662_ (.A1(_1048_),
    .A2(_1072_),
    .B1(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__xor2_1 _3663_ (.A(net299),
    .B(net317),
    .X(_1075_));
 sky130_fd_sc_hd__and2_1 _3664_ (.A(net309),
    .B(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__nor2_1 _3665_ (.A(net309),
    .B(_1075_),
    .Y(_1077_));
 sky130_fd_sc_hd__nor2_1 _3666_ (.A(_1076_),
    .B(_1077_),
    .Y(_1078_));
 sky130_fd_sc_hd__or2_1 _3667_ (.A(net293),
    .B(net312),
    .X(_1079_));
 sky130_fd_sc_hd__nand2_1 _3668_ (.A(net293),
    .B(net312),
    .Y(_1080_));
 sky130_fd_sc_hd__nand3_1 _3669_ (.A(net303),
    .B(_1079_),
    .C(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__a21o_1 _3670_ (.A1(_1079_),
    .A2(_1080_),
    .B1(net303),
    .X(_1082_));
 sky130_fd_sc_hd__nand2_1 _3671_ (.A(_1081_),
    .B(_1082_),
    .Y(_1083_));
 sky130_fd_sc_hd__xor2_1 _3672_ (.A(net296),
    .B(net313),
    .X(_1084_));
 sky130_fd_sc_hd__and2_1 _3673_ (.A(net305),
    .B(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__nor2_1 _3674_ (.A(net306),
    .B(_1084_),
    .Y(_1086_));
 sky130_fd_sc_hd__or2_1 _3675_ (.A(_1085_),
    .B(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__nor2_1 _3676_ (.A(_1083_),
    .B(_1087_),
    .Y(_1088_));
 sky130_fd_sc_hd__or2_1 _3677_ (.A(net297),
    .B(net316),
    .X(_1089_));
 sky130_fd_sc_hd__nand2_1 _3678_ (.A(net297),
    .B(net315),
    .Y(_1090_));
 sky130_fd_sc_hd__a21oi_1 _3679_ (.A1(_1089_),
    .A2(_1090_),
    .B1(net307),
    .Y(_1091_));
 sky130_fd_sc_hd__and3_1 _3680_ (.A(net307),
    .B(_1089_),
    .C(_1090_),
    .X(_1092_));
 sky130_fd_sc_hd__nor2_1 _3681_ (.A(_1091_),
    .B(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__and3_1 _3682_ (.A(_1078_),
    .B(_1088_),
    .C(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__o21bai_1 _3683_ (.A1(_1076_),
    .A2(_1092_),
    .B1_N(_1091_),
    .Y(_1095_));
 sky130_fd_sc_hd__inv_2 _3684_ (.A(_1095_),
    .Y(_1096_));
 sky130_fd_sc_hd__inv_2 _3685_ (.A(_1081_),
    .Y(_1097_));
 sky130_fd_sc_hd__a221o_1 _3686_ (.A1(_1082_),
    .A2(_1085_),
    .B1(_1088_),
    .B2(_1096_),
    .C1(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__a21o_1 _3687_ (.A1(_1074_),
    .A2(_1094_),
    .B1(_1098_),
    .X(_1099_));
 sky130_fd_sc_hd__xor2_1 _3688_ (.A(net291),
    .B(net310),
    .X(_1100_));
 sky130_fd_sc_hd__nand2_1 _3689_ (.A(net301),
    .B(_1100_),
    .Y(_1101_));
 sky130_fd_sc_hd__or2_1 _3690_ (.A(net301),
    .B(_1100_),
    .X(_1102_));
 sky130_fd_sc_hd__nand2_1 _3691_ (.A(_1101_),
    .B(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__or2_1 _3692_ (.A(net289),
    .B(net308),
    .X(_1104_));
 sky130_fd_sc_hd__nand2_1 _3693_ (.A(net289),
    .B(net308),
    .Y(_1105_));
 sky130_fd_sc_hd__a21oi_1 _3694_ (.A1(_1104_),
    .A2(_1105_),
    .B1(net299),
    .Y(_1106_));
 sky130_fd_sc_hd__nand3_1 _3695_ (.A(net300),
    .B(_1104_),
    .C(_1105_),
    .Y(_1107_));
 sky130_fd_sc_hd__or2b_1 _3696_ (.A(_1106_),
    .B_N(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__nor2_1 _3697_ (.A(_1103_),
    .B(_1108_),
    .Y(_1109_));
 sky130_fd_sc_hd__a21oi_1 _3698_ (.A1(_1101_),
    .A2(_1107_),
    .B1(_1106_),
    .Y(_1110_));
 sky130_fd_sc_hd__nand3_1 _3699_ (.A(net298),
    .B(_1040_),
    .C(_1041_),
    .Y(_1111_));
 sky130_fd_sc_hd__nand2_1 _3700_ (.A(_1043_),
    .B(_1111_),
    .Y(_1112_));
 sky130_fd_sc_hd__a211o_1 _3701_ (.A1(_1099_),
    .A2(_1109_),
    .B1(_1110_),
    .C1(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__xor2_1 _3702_ (.A(net282),
    .B(net302),
    .X(_1114_));
 sky130_fd_sc_hd__nand2_1 _3703_ (.A(net293),
    .B(_1114_),
    .Y(_1115_));
 sky130_fd_sc_hd__or2_1 _3704_ (.A(net294),
    .B(_1114_),
    .X(_1116_));
 sky130_fd_sc_hd__nand2_1 _3705_ (.A(_1115_),
    .B(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__or2_1 _3706_ (.A(net280),
    .B(net299),
    .X(_1118_));
 sky130_fd_sc_hd__nand2_1 _3707_ (.A(net280),
    .B(net299),
    .Y(_1119_));
 sky130_fd_sc_hd__nand3_1 _3708_ (.A(net292),
    .B(_1118_),
    .C(_1119_),
    .Y(_1120_));
 sky130_fd_sc_hd__a21oi_1 _3709_ (.A1(_1118_),
    .A2(_1119_),
    .B1(net291),
    .Y(_1121_));
 sky130_fd_sc_hd__inv_2 _3710_ (.A(_1121_),
    .Y(_1122_));
 sky130_fd_sc_hd__nand2_1 _3711_ (.A(_1120_),
    .B(_1122_),
    .Y(_1123_));
 sky130_fd_sc_hd__nor2_1 _3712_ (.A(_1117_),
    .B(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hd__o21ai_1 _3713_ (.A1(_1121_),
    .A2(_1115_),
    .B1(_1120_),
    .Y(_1125_));
 sky130_fd_sc_hd__a31o_1 _3714_ (.A1(_1045_),
    .A2(_1113_),
    .A3(_1124_),
    .B1(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__a21oi_1 _3715_ (.A1(_1033_),
    .A2(_1034_),
    .B1(net289),
    .Y(_1127_));
 sky130_fd_sc_hd__nand3_1 _3716_ (.A(net286),
    .B(_1029_),
    .C(_1030_),
    .Y(_1128_));
 sky130_fd_sc_hd__o21ai_1 _3717_ (.A1(_1031_),
    .A2(_1127_),
    .B1(_1128_),
    .Y(_1129_));
 sky130_fd_sc_hd__or2_1 _3718_ (.A(net284),
    .B(_1022_),
    .X(_1130_));
 sky130_fd_sc_hd__nand2_1 _3719_ (.A(_1023_),
    .B(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__or2b_1 _3720_ (.A(_1027_),
    .B_N(_1026_),
    .X(_1132_));
 sky130_fd_sc_hd__nor2_1 _3721_ (.A(_1131_),
    .B(_1132_),
    .Y(_1133_));
 sky130_fd_sc_hd__o211a_1 _3722_ (.A1(_1036_),
    .A2(_1126_),
    .B1(_1129_),
    .C1(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__a21oi_1 _3723_ (.A1(_1017_),
    .A2(_1018_),
    .B1(net280),
    .Y(_1135_));
 sky130_fd_sc_hd__o21ai_1 _3724_ (.A1(_1020_),
    .A2(_1135_),
    .B1(_1016_),
    .Y(_1136_));
 sky130_fd_sc_hd__o31a_1 _3725_ (.A1(_1021_),
    .A2(_1028_),
    .A3(_1134_),
    .B1(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__and3_1 _3726_ (.A(net276),
    .B(_1011_),
    .C(_1012_),
    .X(_1138_));
 sky130_fd_sc_hd__a21oi_1 _3727_ (.A1(_1013_),
    .A2(_1137_),
    .B1(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__a21oi_1 _3728_ (.A1(_1008_),
    .A2(_1009_),
    .B1(net273),
    .Y(_1140_));
 sky130_fd_sc_hd__or2_1 _3729_ (.A(net272),
    .B(_1006_),
    .X(_1141_));
 sky130_fd_sc_hd__nand2_1 _3730_ (.A(_1007_),
    .B(_1141_),
    .Y(_1142_));
 sky130_fd_sc_hd__a211o_1 _3731_ (.A1(_1010_),
    .A2(_1139_),
    .B1(_1140_),
    .C1(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__nand2_1 _3732_ (.A(_1007_),
    .B(_1143_),
    .Y(_1144_));
 sky130_fd_sc_hd__xnor2_1 _3733_ (.A(_1005_),
    .B(_1144_),
    .Y(_1145_));
 sky130_fd_sc_hd__xnor2_1 _3734_ (.A(_0657_),
    .B(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__nor2_1 _3735_ (.A(_1028_),
    .B(_1134_),
    .Y(_1147_));
 sky130_fd_sc_hd__o21ai_1 _3736_ (.A1(_1147_),
    .A2(_1135_),
    .B1(_1019_),
    .Y(_1148_));
 sky130_fd_sc_hd__inv_2 _3737_ (.A(_1016_),
    .Y(_1149_));
 sky130_fd_sc_hd__nor2_1 _3738_ (.A(_1149_),
    .B(_1020_),
    .Y(_1150_));
 sky130_fd_sc_hd__xnor2_1 _3739_ (.A(_0641_),
    .B(_1150_),
    .Y(_1151_));
 sky130_fd_sc_hd__xor2_1 _3740_ (.A(_1148_),
    .B(_1151_),
    .X(_1152_));
 sky130_fd_sc_hd__nor2_2 _3741_ (.A(_0869_),
    .B(_0998_),
    .Y(_1153_));
 sky130_fd_sc_hd__nand2_2 _3742_ (.A(net265),
    .B(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__clkbuf_2 _3743_ (.A(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__clkbuf_2 _3744_ (.A(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__a21bo_1 _3745_ (.A1(_1099_),
    .A2(_1102_),
    .B1_N(_1101_),
    .X(_1157_));
 sky130_fd_sc_hd__xnor2_1 _3746_ (.A(_1108_),
    .B(_1157_),
    .Y(_1158_));
 sky130_fd_sc_hd__xnor2_1 _3747_ (.A(_0600_),
    .B(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__and2_1 _3748_ (.A(_1156_),
    .B(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__inv_2 _3749_ (.A(_1087_),
    .Y(_1161_));
 sky130_fd_sc_hd__a31o_1 _3750_ (.A1(_1074_),
    .A2(_1078_),
    .A3(_1093_),
    .B1(_1096_),
    .X(_1162_));
 sky130_fd_sc_hd__a21o_1 _3751_ (.A1(_1161_),
    .A2(_1162_),
    .B1(_1085_),
    .X(_1163_));
 sky130_fd_sc_hd__xnor2_2 _3752_ (.A(_1083_),
    .B(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__xnor2_2 _3753_ (.A(_0591_),
    .B(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__xnor2_1 _3754_ (.A(_1087_),
    .B(_1162_),
    .Y(_1166_));
 sky130_fd_sc_hd__xnor2_1 _3755_ (.A(_0524_),
    .B(_1166_),
    .Y(_1167_));
 sky130_fd_sc_hd__a21oi_1 _3756_ (.A1(_1074_),
    .A2(_1078_),
    .B1(_1076_),
    .Y(_1168_));
 sky130_fd_sc_hd__xnor2_2 _3757_ (.A(_1093_),
    .B(_1168_),
    .Y(_1169_));
 sky130_fd_sc_hd__xnor2_2 _3758_ (.A(_0528_),
    .B(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__xor2_1 _3759_ (.A(_1074_),
    .B(_1078_),
    .X(_1171_));
 sky130_fd_sc_hd__xnor2_1 _3760_ (.A(_0586_),
    .B(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__or2b_1 _3761_ (.A(_1073_),
    .B_N(_1048_),
    .X(_1173_));
 sky130_fd_sc_hd__xnor2_2 _3762_ (.A(_1173_),
    .B(_1072_),
    .Y(_1174_));
 sky130_fd_sc_hd__xnor2_1 _3763_ (.A(_0581_),
    .B(_1174_),
    .Y(_1175_));
 sky130_fd_sc_hd__or2b_1 _3764_ (.A(_1071_),
    .B_N(_1051_),
    .X(_1176_));
 sky130_fd_sc_hd__xnor2_2 _3765_ (.A(_1176_),
    .B(_1070_),
    .Y(_1177_));
 sky130_fd_sc_hd__xnor2_2 _3766_ (.A(_0575_),
    .B(_1177_),
    .Y(_1178_));
 sky130_fd_sc_hd__and2b_1 _3767_ (.A_N(_1062_),
    .B(_1060_),
    .X(_1179_));
 sky130_fd_sc_hd__a21oi_1 _3768_ (.A1(net317),
    .A2(_1061_),
    .B1(_1179_),
    .Y(_1180_));
 sky130_fd_sc_hd__xor2_2 _3769_ (.A(_1180_),
    .B(_1067_),
    .X(_1181_));
 sky130_fd_sc_hd__xnor2_1 _3770_ (.A(_0540_),
    .B(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hd__and2b_1 _3771_ (.A_N(_1060_),
    .B(_1062_),
    .X(_1183_));
 sky130_fd_sc_hd__nor2_1 _3772_ (.A(_1179_),
    .B(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__xnor2_1 _3773_ (.A(_0534_),
    .B(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__nand2_1 _3774_ (.A(_1059_),
    .B(_1052_),
    .Y(_1186_));
 sky130_fd_sc_hd__xnor2_2 _3775_ (.A(_1186_),
    .B(_1058_),
    .Y(_1187_));
 sky130_fd_sc_hd__xnor2_1 _3776_ (.A(_0547_),
    .B(_1187_),
    .Y(_1188_));
 sky130_fd_sc_hd__nand2_1 _3777_ (.A(_1057_),
    .B(_1056_),
    .Y(_1189_));
 sky130_fd_sc_hd__xor2_2 _3778_ (.A(_1055_),
    .B(_1189_),
    .X(_1190_));
 sky130_fd_sc_hd__xnor2_1 _3779_ (.A(_0565_),
    .B(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__nand2_1 _3780_ (.A(net315),
    .B(net322),
    .Y(_1192_));
 sky130_fd_sc_hd__xnor2_2 _3781_ (.A(_1053_),
    .B(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__nand3_1 _3782_ (.A(_0557_),
    .B(_0559_),
    .C(_1193_),
    .Y(_1194_));
 sky130_fd_sc_hd__a21o_1 _3783_ (.A1(_0557_),
    .A2(_0559_),
    .B1(_1193_),
    .X(_1195_));
 sky130_fd_sc_hd__or2_1 _3784_ (.A(net315),
    .B(net322),
    .X(_1196_));
 sky130_fd_sc_hd__nand2_2 _3785_ (.A(_1192_),
    .B(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__xor2_2 _3786_ (.A(_0553_),
    .B(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__a21o_1 _3787_ (.A1(_1194_),
    .A2(_1195_),
    .B1(_1198_),
    .X(_1199_));
 sky130_fd_sc_hd__or3_1 _3788_ (.A(_1188_),
    .B(_1191_),
    .C(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__or3_1 _3789_ (.A(_1182_),
    .B(_1185_),
    .C(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__or4_1 _3790_ (.A(_1172_),
    .B(_1175_),
    .C(_1178_),
    .D(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__or3_1 _3791_ (.A(_1167_),
    .B(_1170_),
    .C(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__xnor2_1 _3792_ (.A(_1099_),
    .B(_1103_),
    .Y(_1204_));
 sky130_fd_sc_hd__xnor2_2 _3793_ (.A(_0606_),
    .B(_1204_),
    .Y(_1205_));
 sky130_fd_sc_hd__o31a_1 _3794_ (.A1(_1165_),
    .A2(_1203_),
    .A3(_1205_),
    .B1(_1156_),
    .X(_1206_));
 sky130_fd_sc_hd__a21o_1 _3795_ (.A1(_1099_),
    .A2(_1109_),
    .B1(_1110_),
    .X(_1207_));
 sky130_fd_sc_hd__nand2_1 _3796_ (.A(_1042_),
    .B(_1111_),
    .Y(_1208_));
 sky130_fd_sc_hd__xnor2_1 _3797_ (.A(_1207_),
    .B(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__xnor2_1 _3798_ (.A(_0611_),
    .B(_1209_),
    .Y(_1210_));
 sky130_fd_sc_hd__nor2_1 _3799_ (.A(_1000_),
    .B(_1210_),
    .Y(_1211_));
 sky130_fd_sc_hd__or3_1 _3800_ (.A(_1160_),
    .B(_1206_),
    .C(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__nand2_1 _3801_ (.A(_1045_),
    .B(_1113_),
    .Y(_1213_));
 sky130_fd_sc_hd__xor2_2 _3802_ (.A(_1213_),
    .B(_1117_),
    .X(_1214_));
 sky130_fd_sc_hd__xor2_1 _3803_ (.A(_0616_),
    .B(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__o21ai_1 _3804_ (.A1(_1213_),
    .A2(_1117_),
    .B1(_1115_),
    .Y(_1216_));
 sky130_fd_sc_hd__xor2_1 _3805_ (.A(_0619_),
    .B(_1123_),
    .X(_1217_));
 sky130_fd_sc_hd__xnor2_2 _3806_ (.A(_1216_),
    .B(_1217_),
    .Y(_1218_));
 sky130_fd_sc_hd__nand2_1 _3807_ (.A(_1039_),
    .B(_1043_),
    .Y(_1219_));
 sky130_fd_sc_hd__a21bo_1 _3808_ (.A1(_1042_),
    .A2(_1207_),
    .B1_N(_1111_),
    .X(_1220_));
 sky130_fd_sc_hd__xnor2_1 _3809_ (.A(_1219_),
    .B(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__xnor2_2 _3810_ (.A(_0501_),
    .B(_1221_),
    .Y(_1222_));
 sky130_fd_sc_hd__nand2_1 _3811_ (.A(_1156_),
    .B(_1222_),
    .Y(_1223_));
 sky130_fd_sc_hd__and4b_2 _3812_ (.A_N(_1212_),
    .B(_1215_),
    .C(_1218_),
    .D(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__nor2_1 _3813_ (.A(_1035_),
    .B(_1127_),
    .Y(_1225_));
 sky130_fd_sc_hd__xnor2_1 _3814_ (.A(_1126_),
    .B(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__xor2_2 _3815_ (.A(_0624_),
    .B(_1226_),
    .X(_1227_));
 sky130_fd_sc_hd__inv_2 _3816_ (.A(_1227_),
    .Y(_1228_));
 sky130_fd_sc_hd__nand2_1 _3817_ (.A(_1128_),
    .B(_1032_),
    .Y(_1229_));
 sky130_fd_sc_hd__a21oi_1 _3818_ (.A1(_1126_),
    .A2(_1225_),
    .B1(_1035_),
    .Y(_1230_));
 sky130_fd_sc_hd__xnor2_2 _3819_ (.A(_1229_),
    .B(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__xor2_4 _3820_ (.A(_0496_),
    .B(_1231_),
    .X(_1232_));
 sky130_fd_sc_hd__nor2_1 _3821_ (.A(_1228_),
    .B(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__o21ai_1 _3822_ (.A1(_1036_),
    .A2(_1126_),
    .B1(_1129_),
    .Y(_1234_));
 sky130_fd_sc_hd__or2_1 _3823_ (.A(_1234_),
    .B(_1131_),
    .X(_1235_));
 sky130_fd_sc_hd__nand2_1 _3824_ (.A(_1234_),
    .B(_1131_),
    .Y(_1236_));
 sky130_fd_sc_hd__nand2_1 _3825_ (.A(_1235_),
    .B(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__xnor2_2 _3826_ (.A(_0629_),
    .B(_1237_),
    .Y(_1238_));
 sky130_fd_sc_hd__nand2_1 _3827_ (.A(_1023_),
    .B(_1235_),
    .Y(_1239_));
 sky130_fd_sc_hd__xor2_1 _3828_ (.A(_0486_),
    .B(_1132_),
    .X(_1240_));
 sky130_fd_sc_hd__xnor2_1 _3829_ (.A(_1239_),
    .B(_1240_),
    .Y(_1241_));
 sky130_fd_sc_hd__a41o_1 _3830_ (.A1(_1224_),
    .A2(_1233_),
    .A3(_1238_),
    .A4(_1241_),
    .B1(_1000_),
    .X(_1242_));
 sky130_fd_sc_hd__clkbuf_2 _3831_ (.A(_1156_),
    .X(_1243_));
 sky130_fd_sc_hd__inv_2 _3832_ (.A(_1135_),
    .Y(_1244_));
 sky130_fd_sc_hd__nand2_1 _3833_ (.A(_1019_),
    .B(_1244_),
    .Y(_1245_));
 sky130_fd_sc_hd__xnor2_1 _3834_ (.A(_1147_),
    .B(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__xor2_2 _3835_ (.A(_0635_),
    .B(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__nand2_1 _3836_ (.A(_1243_),
    .B(_1247_),
    .Y(_1248_));
 sky130_fd_sc_hd__nand3b_2 _3837_ (.A_N(_1152_),
    .B(_1242_),
    .C(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__inv_2 _3838_ (.A(_1140_),
    .Y(_1250_));
 sky130_fd_sc_hd__nand2_1 _3839_ (.A(_1010_),
    .B(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__xor2_1 _3840_ (.A(_1139_),
    .B(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__and3_1 _3841_ (.A(_0474_),
    .B(_0475_),
    .C(_1252_),
    .X(_1253_));
 sky130_fd_sc_hd__a21oi_1 _3842_ (.A1(_0474_),
    .A2(_0475_),
    .B1(_1252_),
    .Y(_1254_));
 sky130_fd_sc_hd__or2b_1 _3843_ (.A(_1138_),
    .B_N(_1013_),
    .X(_1255_));
 sky130_fd_sc_hd__xnor2_1 _3844_ (.A(_1255_),
    .B(_1137_),
    .Y(_1256_));
 sky130_fd_sc_hd__xnor2_2 _3845_ (.A(_0647_),
    .B(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__o21ai_1 _3846_ (.A1(_1253_),
    .A2(_1254_),
    .B1(_1257_),
    .Y(_1258_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3847_ (.A(_1243_),
    .X(_1259_));
 sky130_fd_sc_hd__o21ai_1 _3848_ (.A1(_1249_),
    .A2(_1258_),
    .B1(_1259_),
    .Y(_1260_));
 sky130_fd_sc_hd__a21oi_1 _3849_ (.A1(_1010_),
    .A2(_1139_),
    .B1(_1140_),
    .Y(_1261_));
 sky130_fd_sc_hd__xnor2_1 _3850_ (.A(_1142_),
    .B(_1261_),
    .Y(_1262_));
 sky130_fd_sc_hd__xnor2_2 _3851_ (.A(_0652_),
    .B(_1262_),
    .Y(_1263_));
 sky130_fd_sc_hd__nand2_1 _3852_ (.A(_1259_),
    .B(_1263_),
    .Y(_1264_));
 sky130_fd_sc_hd__and3b_1 _3853_ (.A_N(_1146_),
    .B(_1260_),
    .C(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__nand2_1 _3854_ (.A(net268),
    .B(net276),
    .Y(_1266_));
 sky130_fd_sc_hd__or2_1 _3855_ (.A(net268),
    .B(net276),
    .X(_1267_));
 sky130_fd_sc_hd__nand2_1 _3856_ (.A(_1266_),
    .B(_1267_),
    .Y(_1268_));
 sky130_fd_sc_hd__nor2_1 _3857_ (.A(net270),
    .B(net279),
    .Y(_1269_));
 sky130_fd_sc_hd__a31o_1 _3858_ (.A1(_1007_),
    .A2(_1143_),
    .A3(_1003_),
    .B1(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__xor2_1 _3859_ (.A(_1268_),
    .B(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__xnor2_2 _3860_ (.A(_0665_),
    .B(_1271_),
    .Y(_1272_));
 sky130_fd_sc_hd__nand2_1 _3861_ (.A(_1259_),
    .B(_1272_),
    .Y(_1273_));
 sky130_fd_sc_hd__o21a_1 _3862_ (.A1(_1268_),
    .A2(_1270_),
    .B1(_1266_),
    .X(_1274_));
 sky130_fd_sc_hd__nor2_1 _3863_ (.A(net267),
    .B(net274),
    .Y(_1275_));
 sky130_fd_sc_hd__and2_1 _3864_ (.A(net267),
    .B(net273),
    .X(_1276_));
 sky130_fd_sc_hd__or2_1 _3865_ (.A(_1275_),
    .B(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__xnor2_1 _3866_ (.A(_1274_),
    .B(_1277_),
    .Y(_1278_));
 sky130_fd_sc_hd__xnor2_1 _3867_ (.A(_2161_),
    .B(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__o211a_1 _3868_ (.A1(_1002_),
    .A2(_1265_),
    .B1(_1273_),
    .C1(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__nor2_1 _3869_ (.A(_1002_),
    .B(_1280_),
    .Y(_1281_));
 sky130_fd_sc_hd__nand2_1 _3870_ (.A(net266),
    .B(net272),
    .Y(_1282_));
 sky130_fd_sc_hd__or2_1 _3871_ (.A(net266),
    .B(net272),
    .X(_1283_));
 sky130_fd_sc_hd__nand2_1 _3872_ (.A(_1282_),
    .B(_1283_),
    .Y(_1284_));
 sky130_fd_sc_hd__o21ba_1 _3873_ (.A1(_1274_),
    .A2(_1275_),
    .B1_N(_1276_),
    .X(_1285_));
 sky130_fd_sc_hd__xor2_1 _3874_ (.A(_1284_),
    .B(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__xnor2_2 _3875_ (.A(_0685_),
    .B(_1286_),
    .Y(_1287_));
 sky130_fd_sc_hd__xnor2_1 _3876_ (.A(_1281_),
    .B(_1287_),
    .Y(_1288_));
 sky130_fd_sc_hd__nand2_1 _3877_ (.A(net323),
    .B(_1288_),
    .Y(_1289_));
 sky130_fd_sc_hd__or2_1 _3878_ (.A(_1002_),
    .B(_1265_),
    .X(_1290_));
 sky130_fd_sc_hd__xnor2_1 _3879_ (.A(_1272_),
    .B(_1290_),
    .Y(_1291_));
 sky130_fd_sc_hd__nand2_1 _3880_ (.A(net325),
    .B(_1291_),
    .Y(_1292_));
 sky130_fd_sc_hd__xor2_1 _3881_ (.A(_1222_),
    .B(_1212_),
    .X(_1293_));
 sky130_fd_sc_hd__nand2_1 _3882_ (.A(net350),
    .B(_1293_),
    .Y(_1294_));
 sky130_fd_sc_hd__or2_1 _3883_ (.A(_1160_),
    .B(_1206_),
    .X(_1295_));
 sky130_fd_sc_hd__xnor2_1 _3884_ (.A(_1295_),
    .B(_1210_),
    .Y(_1296_));
 sky130_fd_sc_hd__and2_1 _3885_ (.A(net353),
    .B(_1296_),
    .X(_1297_));
 sky130_fd_sc_hd__xor2_1 _3886_ (.A(_1159_),
    .B(_1206_),
    .X(_1298_));
 sky130_fd_sc_hd__or2_1 _3887_ (.A(net355),
    .B(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__inv_2 _3888_ (.A(_1299_),
    .Y(_1300_));
 sky130_fd_sc_hd__o21ai_1 _3889_ (.A1(_1165_),
    .A2(_1203_),
    .B1(_1243_),
    .Y(_1301_));
 sky130_fd_sc_hd__xnor2_1 _3890_ (.A(_1301_),
    .B(_1205_),
    .Y(_1302_));
 sky130_fd_sc_hd__nand2_1 _3891_ (.A(net356),
    .B(_1302_),
    .Y(_1303_));
 sky130_fd_sc_hd__and2_1 _3892_ (.A(net354),
    .B(_1298_),
    .X(_1304_));
 sky130_fd_sc_hd__o21ba_1 _3893_ (.A1(_1300_),
    .A2(_1303_),
    .B1_N(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__or2_1 _3894_ (.A(net356),
    .B(_1302_),
    .X(_1306_));
 sky130_fd_sc_hd__nand2_1 _3895_ (.A(_1303_),
    .B(_1306_),
    .Y(_1307_));
 sky130_fd_sc_hd__and2_1 _3896_ (.A(_1243_),
    .B(_1203_),
    .X(_1308_));
 sky130_fd_sc_hd__xor2_1 _3897_ (.A(_1165_),
    .B(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__nor2_1 _3898_ (.A(net358),
    .B(_1309_),
    .Y(_1310_));
 sky130_fd_sc_hd__nand2_1 _3899_ (.A(_1155_),
    .B(_1202_),
    .Y(_1311_));
 sky130_fd_sc_hd__xnor2_1 _3900_ (.A(_1170_),
    .B(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hd__nor2_1 _3901_ (.A(net362),
    .B(_1312_),
    .Y(_1313_));
 sky130_fd_sc_hd__o31a_1 _3902_ (.A1(_1175_),
    .A2(_1178_),
    .A3(_1201_),
    .B1(_1155_),
    .X(_1314_));
 sky130_fd_sc_hd__xor2_1 _3903_ (.A(_1172_),
    .B(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__nand2_1 _3904_ (.A(net364),
    .B(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__or2_1 _3905_ (.A(net364),
    .B(_1315_),
    .X(_1317_));
 sky130_fd_sc_hd__and2_1 _3906_ (.A(_1316_),
    .B(_1317_),
    .X(_1318_));
 sky130_fd_sc_hd__inv_2 _3907_ (.A(_1318_),
    .Y(_1319_));
 sky130_fd_sc_hd__o21ai_1 _3908_ (.A1(_1178_),
    .A2(_1201_),
    .B1(_1156_),
    .Y(_1320_));
 sky130_fd_sc_hd__xnor2_1 _3909_ (.A(_1175_),
    .B(_1320_),
    .Y(_1321_));
 sky130_fd_sc_hd__or2_1 _3910_ (.A(net366),
    .B(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__nand2_1 _3911_ (.A(_1155_),
    .B(_1201_),
    .Y(_1323_));
 sky130_fd_sc_hd__xnor2_1 _3912_ (.A(_1178_),
    .B(_1323_),
    .Y(_1324_));
 sky130_fd_sc_hd__xor2_1 _3913_ (.A(net368),
    .B(_1324_),
    .X(_1325_));
 sky130_fd_sc_hd__o21a_1 _3914_ (.A1(_1191_),
    .A2(_1199_),
    .B1(_1154_),
    .X(_1326_));
 sky130_fd_sc_hd__a21o_1 _3915_ (.A1(_1155_),
    .A2(_1188_),
    .B1(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__a21oi_1 _3916_ (.A1(_1155_),
    .A2(_1185_),
    .B1(_1327_),
    .Y(_1328_));
 sky130_fd_sc_hd__xnor2_1 _3917_ (.A(_1182_),
    .B(_1328_),
    .Y(_1329_));
 sky130_fd_sc_hd__xor2_1 _3918_ (.A(net371),
    .B(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__xor2_1 _3919_ (.A(_1188_),
    .B(_1326_),
    .X(_1331_));
 sky130_fd_sc_hd__xor2_1 _3920_ (.A(net373),
    .B(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__a22o_1 _3921_ (.A1(_1154_),
    .A2(_1198_),
    .B1(_1194_),
    .B2(_1195_),
    .X(_1333_));
 sky130_fd_sc_hd__nand4_1 _3922_ (.A(_1154_),
    .B(_1198_),
    .C(_1194_),
    .D(_1195_),
    .Y(_1334_));
 sky130_fd_sc_hd__a21o_1 _3923_ (.A1(_1333_),
    .A2(_1334_),
    .B1(\workunit1[1] ),
    .X(_1335_));
 sky130_fd_sc_hd__and3_1 _3924_ (.A(\workunit1[1] ),
    .B(_1333_),
    .C(_1334_),
    .X(_1336_));
 sky130_fd_sc_hd__a31o_1 _3925_ (.A1(net376),
    .A2(_1198_),
    .A3(_1335_),
    .B1(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__nand3_1 _3926_ (.A(_1154_),
    .B(_1191_),
    .C(_1199_),
    .Y(_1338_));
 sky130_fd_sc_hd__a21o_1 _3927_ (.A1(_1154_),
    .A2(_1199_),
    .B1(_1191_),
    .X(_1339_));
 sky130_fd_sc_hd__a21o_1 _3928_ (.A1(_1338_),
    .A2(_1339_),
    .B1(net374),
    .X(_1340_));
 sky130_fd_sc_hd__and3_1 _3929_ (.A(net374),
    .B(_1338_),
    .C(_1339_),
    .X(_1341_));
 sky130_fd_sc_hd__a21o_1 _3930_ (.A1(_1337_),
    .A2(_1340_),
    .B1(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__and2_1 _3931_ (.A(net373),
    .B(_1331_),
    .X(_1343_));
 sky130_fd_sc_hd__a21o_1 _3932_ (.A1(_1332_),
    .A2(_1342_),
    .B1(_1343_),
    .X(_1344_));
 sky130_fd_sc_hd__xor2_1 _3933_ (.A(_1185_),
    .B(_1327_),
    .X(_1345_));
 sky130_fd_sc_hd__xor2_1 _3934_ (.A(net372),
    .B(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__and2_1 _3935_ (.A(net372),
    .B(_1345_),
    .X(_1347_));
 sky130_fd_sc_hd__a21o_1 _3936_ (.A1(_1344_),
    .A2(_1346_),
    .B1(_1347_),
    .X(_1348_));
 sky130_fd_sc_hd__and2_1 _3937_ (.A(net371),
    .B(_1329_),
    .X(_1349_));
 sky130_fd_sc_hd__a21o_1 _3938_ (.A1(_1330_),
    .A2(_1348_),
    .B1(_1349_),
    .X(_1350_));
 sky130_fd_sc_hd__and2_1 _3939_ (.A(net368),
    .B(_1324_),
    .X(_1351_));
 sky130_fd_sc_hd__a21o_1 _3940_ (.A1(_1325_),
    .A2(_1350_),
    .B1(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__and2_1 _3941_ (.A(net366),
    .B(_1321_),
    .X(_1353_));
 sky130_fd_sc_hd__a21oi_1 _3942_ (.A1(_1322_),
    .A2(_1352_),
    .B1(_1353_),
    .Y(_1354_));
 sky130_fd_sc_hd__and2_1 _3943_ (.A(net362),
    .B(_1312_),
    .X(_1355_));
 sky130_fd_sc_hd__inv_2 _3944_ (.A(_1355_),
    .Y(_1356_));
 sky130_fd_sc_hd__o211a_1 _3945_ (.A1(_1319_),
    .A2(_1354_),
    .B1(_1356_),
    .C1(_1316_),
    .X(_1357_));
 sky130_fd_sc_hd__o21ai_1 _3946_ (.A1(_1170_),
    .A2(_1202_),
    .B1(_1156_),
    .Y(_1358_));
 sky130_fd_sc_hd__xnor2_1 _3947_ (.A(_1167_),
    .B(_1358_),
    .Y(_1359_));
 sky130_fd_sc_hd__nand2_1 _3948_ (.A(net360),
    .B(_1359_),
    .Y(_1360_));
 sky130_fd_sc_hd__or2_1 _3949_ (.A(net360),
    .B(_1359_),
    .X(_1361_));
 sky130_fd_sc_hd__and2_1 _3950_ (.A(_1360_),
    .B(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__inv_2 _3951_ (.A(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__nand2_1 _3952_ (.A(net358),
    .B(_1309_),
    .Y(_1364_));
 sky130_fd_sc_hd__o311a_1 _3953_ (.A1(_1313_),
    .A2(_1357_),
    .A3(_1363_),
    .B1(_1360_),
    .C1(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__or2_1 _3954_ (.A(_1304_),
    .B(_1300_),
    .X(_1366_));
 sky130_fd_sc_hd__or4_1 _3955_ (.A(_1307_),
    .B(_1310_),
    .C(_1365_),
    .D(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__nor2_1 _3956_ (.A(net353),
    .B(_1296_),
    .Y(_1368_));
 sky130_fd_sc_hd__nor2_1 _3957_ (.A(_1297_),
    .B(_1368_),
    .Y(_1369_));
 sky130_fd_sc_hd__inv_2 _3958_ (.A(_1369_),
    .Y(_1370_));
 sky130_fd_sc_hd__a21oi_1 _3959_ (.A1(_1305_),
    .A2(_1367_),
    .B1(_1370_),
    .Y(_1371_));
 sky130_fd_sc_hd__or2_1 _3960_ (.A(net350),
    .B(_1293_),
    .X(_1372_));
 sky130_fd_sc_hd__and2_1 _3961_ (.A(_1294_),
    .B(_1372_),
    .X(_1373_));
 sky130_fd_sc_hd__o21ai_2 _3962_ (.A1(_1297_),
    .A2(_1371_),
    .B1(_1373_),
    .Y(_1374_));
 sky130_fd_sc_hd__a21o_1 _3963_ (.A1(_1224_),
    .A2(_1227_),
    .B1(_1001_),
    .X(_1375_));
 sky130_fd_sc_hd__xnor2_2 _3964_ (.A(_1232_),
    .B(_1375_),
    .Y(_1376_));
 sky130_fd_sc_hd__xnor2_1 _3965_ (.A(net341),
    .B(_1376_),
    .Y(_1377_));
 sky130_fd_sc_hd__or3_1 _3966_ (.A(_1000_),
    .B(_1224_),
    .C(_1228_),
    .X(_1378_));
 sky130_fd_sc_hd__o21ai_1 _3967_ (.A1(_1001_),
    .A2(_1224_),
    .B1(_1228_),
    .Y(_1379_));
 sky130_fd_sc_hd__a21boi_1 _3968_ (.A1(_1378_),
    .A2(_1379_),
    .B1_N(net344),
    .Y(_1380_));
 sky130_fd_sc_hd__and3b_1 _3969_ (.A_N(net344),
    .B(_1378_),
    .C(_1379_),
    .X(_1381_));
 sky130_fd_sc_hd__xnor2_1 _3970_ (.A(_0616_),
    .B(_1214_),
    .Y(_1382_));
 sky130_fd_sc_hd__o31a_1 _3971_ (.A1(_1222_),
    .A2(_1212_),
    .A3(_1382_),
    .B1(_1243_),
    .X(_1383_));
 sky130_fd_sc_hd__xnor2_1 _3972_ (.A(_1218_),
    .B(_1383_),
    .Y(_1384_));
 sky130_fd_sc_hd__nor2_1 _3973_ (.A(net346),
    .B(_1384_),
    .Y(_1385_));
 sky130_fd_sc_hd__or3_1 _3974_ (.A(_1380_),
    .B(_1381_),
    .C(_1385_),
    .X(_1386_));
 sky130_fd_sc_hd__and2_1 _3975_ (.A(net346),
    .B(_1384_),
    .X(_1387_));
 sky130_fd_sc_hd__or2b_1 _3976_ (.A(_1212_),
    .B_N(_1223_),
    .X(_1388_));
 sky130_fd_sc_hd__xnor2_1 _3977_ (.A(_1388_),
    .B(_1215_),
    .Y(_1389_));
 sky130_fd_sc_hd__nor2_1 _3978_ (.A(net348),
    .B(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__and2_1 _3979_ (.A(net348),
    .B(_1389_),
    .X(_1391_));
 sky130_fd_sc_hd__or2_1 _3980_ (.A(_1390_),
    .B(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__or4_1 _3981_ (.A(_1377_),
    .B(_1386_),
    .C(_1387_),
    .D(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__a21bo_1 _3982_ (.A1(_1242_),
    .A2(_1248_),
    .B1_N(_1152_),
    .X(_1394_));
 sky130_fd_sc_hd__nand2_1 _3983_ (.A(_1249_),
    .B(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hd__xnor2_1 _3984_ (.A(net334),
    .B(_1395_),
    .Y(_1396_));
 sky130_fd_sc_hd__xnor2_1 _3985_ (.A(_1242_),
    .B(_1247_),
    .Y(_1397_));
 sky130_fd_sc_hd__xnor2_1 _3986_ (.A(net336),
    .B(_1397_),
    .Y(_1398_));
 sky130_fd_sc_hd__inv_2 _3987_ (.A(_1398_),
    .Y(_1399_));
 sky130_fd_sc_hd__o21ai_1 _3988_ (.A1(_1228_),
    .A2(_1232_),
    .B1(_1243_),
    .Y(_1400_));
 sky130_fd_sc_hd__o211a_1 _3989_ (.A1(_1001_),
    .A2(_1224_),
    .B1(_1400_),
    .C1(_1238_),
    .X(_1401_));
 sky130_fd_sc_hd__a211oi_1 _3990_ (.A1(_1224_),
    .A2(_1233_),
    .B1(_1238_),
    .C1(_1001_),
    .Y(_1402_));
 sky130_fd_sc_hd__nor2_1 _3991_ (.A(_1401_),
    .B(_1402_),
    .Y(_1403_));
 sky130_fd_sc_hd__and2_1 _3992_ (.A(net339),
    .B(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__nor2_1 _3993_ (.A(net339),
    .B(_1403_),
    .Y(_1405_));
 sky130_fd_sc_hd__nor2_1 _3994_ (.A(_1404_),
    .B(_1405_),
    .Y(_1406_));
 sky130_fd_sc_hd__inv_2 _3995_ (.A(\workunit1[21] ),
    .Y(_1407_));
 sky130_fd_sc_hd__or3b_1 _3996_ (.A(_1001_),
    .B(_1401_),
    .C_N(_1241_),
    .X(_1408_));
 sky130_fd_sc_hd__o21bai_2 _3997_ (.A1(_1002_),
    .A2(_1401_),
    .B1_N(_1241_),
    .Y(_1409_));
 sky130_fd_sc_hd__and3_1 _3998_ (.A(_1407_),
    .B(_1408_),
    .C(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__a21oi_1 _3999_ (.A1(_1408_),
    .A2(_1409_),
    .B1(_1407_),
    .Y(_1411_));
 sky130_fd_sc_hd__nor2_1 _4000_ (.A(_1410_),
    .B(_1411_),
    .Y(_1412_));
 sky130_fd_sc_hd__nand4_1 _4001_ (.A(_1396_),
    .B(_1399_),
    .C(_1406_),
    .D(_1412_),
    .Y(_1413_));
 sky130_fd_sc_hd__a211o_1 _4002_ (.A1(_1294_),
    .A2(_1374_),
    .B1(_1393_),
    .C1(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__nor2_1 _4003_ (.A(_1377_),
    .B(_1386_),
    .Y(_1415_));
 sky130_fd_sc_hd__or2_1 _4004_ (.A(_1387_),
    .B(_1391_),
    .X(_1416_));
 sky130_fd_sc_hd__o21a_1 _4005_ (.A1(net341),
    .A2(_1376_),
    .B1(_1380_),
    .X(_1417_));
 sky130_fd_sc_hd__a221oi_1 _4006_ (.A1(net341),
    .A2(_1376_),
    .B1(_1415_),
    .B2(_1416_),
    .C1(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__nand3_2 _4007_ (.A(_1407_),
    .B(_1408_),
    .C(_1409_),
    .Y(_1419_));
 sky130_fd_sc_hd__o2111ai_1 _4008_ (.A1(_1404_),
    .A2(_1411_),
    .B1(_1419_),
    .C1(_1396_),
    .D1(_1399_),
    .Y(_1420_));
 sky130_fd_sc_hd__inv_2 _4009_ (.A(net334),
    .Y(_1421_));
 sky130_fd_sc_hd__nand2_1 _4010_ (.A(_1421_),
    .B(_1395_),
    .Y(_1422_));
 sky130_fd_sc_hd__and2_1 _4011_ (.A(net336),
    .B(_1397_),
    .X(_1423_));
 sky130_fd_sc_hd__nor2_1 _4012_ (.A(_1421_),
    .B(_1395_),
    .Y(_1424_));
 sky130_fd_sc_hd__a21oi_1 _4013_ (.A1(_1422_),
    .A2(_1423_),
    .B1(_1424_),
    .Y(_1425_));
 sky130_fd_sc_hd__o211a_1 _4014_ (.A1(_1413_),
    .A2(_1418_),
    .B1(_1420_),
    .C1(_1425_),
    .X(_1426_));
 sky130_fd_sc_hd__inv_2 _4015_ (.A(_1257_),
    .Y(_1427_));
 sky130_fd_sc_hd__nand2_1 _4016_ (.A(_1259_),
    .B(_1249_),
    .Y(_1428_));
 sky130_fd_sc_hd__xnor2_1 _4017_ (.A(_1427_),
    .B(_1428_),
    .Y(_1429_));
 sky130_fd_sc_hd__and2_1 _4018_ (.A(net333),
    .B(_1429_),
    .X(_1430_));
 sky130_fd_sc_hd__nor2_1 _4019_ (.A(net333),
    .B(_1429_),
    .Y(_1431_));
 sky130_fd_sc_hd__or2_1 _4020_ (.A(_1430_),
    .B(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__nor2_1 _4021_ (.A(_1253_),
    .B(_1254_),
    .Y(_1433_));
 sky130_fd_sc_hd__o21ai_1 _4022_ (.A1(_1249_),
    .A2(_1427_),
    .B1(_1259_),
    .Y(_1434_));
 sky130_fd_sc_hd__xnor2_2 _4023_ (.A(_1433_),
    .B(_1434_),
    .Y(_1435_));
 sky130_fd_sc_hd__xnor2_1 _4024_ (.A(net331),
    .B(_1435_),
    .Y(_1436_));
 sky130_fd_sc_hd__o31ai_1 _4025_ (.A1(_1263_),
    .A2(_1249_),
    .A3(_1258_),
    .B1(_1259_),
    .Y(_1437_));
 sky130_fd_sc_hd__xnor2_1 _4026_ (.A(_1437_),
    .B(_1146_),
    .Y(_1438_));
 sky130_fd_sc_hd__xnor2_1 _4027_ (.A(net326),
    .B(_1438_),
    .Y(_1439_));
 sky130_fd_sc_hd__xnor2_1 _4028_ (.A(_1263_),
    .B(_1260_),
    .Y(_1440_));
 sky130_fd_sc_hd__xnor2_2 _4029_ (.A(net329),
    .B(_1440_),
    .Y(_1441_));
 sky130_fd_sc_hd__or3_1 _4030_ (.A(_1436_),
    .B(_1439_),
    .C(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__a211o_1 _4031_ (.A1(_1414_),
    .A2(_1426_),
    .B1(_1432_),
    .C1(_1442_),
    .X(_1443_));
 sky130_fd_sc_hd__nor2_1 _4032_ (.A(net331),
    .B(_1435_),
    .Y(_1444_));
 sky130_fd_sc_hd__inv_2 _4033_ (.A(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__nor2_1 _4034_ (.A(_1439_),
    .B(_1441_),
    .Y(_1446_));
 sky130_fd_sc_hd__a21o_1 _4035_ (.A1(net331),
    .A2(_1435_),
    .B1(_1430_),
    .X(_1447_));
 sky130_fd_sc_hd__and2_1 _4036_ (.A(net329),
    .B(_1440_),
    .X(_1448_));
 sky130_fd_sc_hd__a21o_1 _4037_ (.A1(net326),
    .A2(_1438_),
    .B1(_1448_),
    .X(_1449_));
 sky130_fd_sc_hd__or2_1 _4038_ (.A(net326),
    .B(_1438_),
    .X(_1450_));
 sky130_fd_sc_hd__a32oi_2 _4039_ (.A1(_1445_),
    .A2(_1446_),
    .A3(_1447_),
    .B1(_1449_),
    .B2(_1450_),
    .Y(_1451_));
 sky130_fd_sc_hd__xnor2_1 _4040_ (.A(net325),
    .B(_1291_),
    .Y(_1452_));
 sky130_fd_sc_hd__a21o_1 _4041_ (.A1(_1443_),
    .A2(_1451_),
    .B1(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__a21oi_1 _4042_ (.A1(_1290_),
    .A2(_1273_),
    .B1(_1279_),
    .Y(_1454_));
 sky130_fd_sc_hd__nor2_1 _4043_ (.A(_1280_),
    .B(_1454_),
    .Y(_1455_));
 sky130_fd_sc_hd__nand2_1 _4044_ (.A(net324),
    .B(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__nor2_1 _4045_ (.A(net324),
    .B(_1455_),
    .Y(_1457_));
 sky130_fd_sc_hd__xnor2_1 _4046_ (.A(net323),
    .B(_1288_),
    .Y(_1458_));
 sky130_fd_sc_hd__a311o_1 _4047_ (.A1(_1292_),
    .A2(_1453_),
    .A3(_1456_),
    .B1(_1457_),
    .C1(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__a21oi_1 _4048_ (.A1(_1280_),
    .A2(_1287_),
    .B1(_1002_),
    .Y(_1460_));
 sky130_fd_sc_hd__o21a_1 _4049_ (.A1(_1284_),
    .A2(_1285_),
    .B1(_1282_),
    .X(_1461_));
 sky130_fd_sc_hd__xor2_1 _4050_ (.A(net270),
    .B(_0858_),
    .X(_1462_));
 sky130_fd_sc_hd__xnor2_1 _4051_ (.A(_1461_),
    .B(_1462_),
    .Y(_1463_));
 sky130_fd_sc_hd__xnor2_1 _4052_ (.A(_0856_),
    .B(_1463_),
    .Y(_1464_));
 sky130_fd_sc_hd__xnor2_1 _4053_ (.A(_1460_),
    .B(_1464_),
    .Y(_1465_));
 sky130_fd_sc_hd__and3_1 _4054_ (.A(_1289_),
    .B(_1459_),
    .C(_1465_),
    .X(_1466_));
 sky130_fd_sc_hd__a21oi_1 _4055_ (.A1(_1289_),
    .A2(_1459_),
    .B1(_1465_),
    .Y(_1467_));
 sky130_fd_sc_hd__buf_2 _4056_ (.A(_1153_),
    .X(_1468_));
 sky130_fd_sc_hd__clkbuf_2 _4057_ (.A(_1468_),
    .X(_1469_));
 sky130_fd_sc_hd__o21ai_1 _4058_ (.A1(_1466_),
    .A2(_1467_),
    .B1(_1469_),
    .Y(_1470_));
 sky130_fd_sc_hd__a21o_1 _4059_ (.A1(net531),
    .A2(_0874_),
    .B1(_1469_),
    .X(_1471_));
 sky130_fd_sc_hd__nor2_1 _4060_ (.A(_0872_),
    .B(_1153_),
    .Y(_1472_));
 sky130_fd_sc_hd__buf_2 _4061_ (.A(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__clkbuf_2 _4062_ (.A(_1473_),
    .X(_1474_));
 sky130_fd_sc_hd__a22o_1 _4063_ (.A1(_1470_),
    .A2(_1471_),
    .B1(_1474_),
    .B2(\workunit1[31] ),
    .X(_0320_));
 sky130_fd_sc_hd__buf_2 _4064_ (.A(_1469_),
    .X(_1475_));
 sky130_fd_sc_hd__a31o_1 _4065_ (.A1(_1292_),
    .A2(_1453_),
    .A3(_1456_),
    .B1(_1457_),
    .X(_1476_));
 sky130_fd_sc_hd__nand2_1 _4066_ (.A(_1458_),
    .B(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__buf_2 _4067_ (.A(_1472_),
    .X(_1478_));
 sky130_fd_sc_hd__a22o_1 _4068_ (.A1(net488),
    .A2(_0874_),
    .B1(_1478_),
    .B2(net323),
    .X(_1479_));
 sky130_fd_sc_hd__a31o_1 _4069_ (.A1(_1475_),
    .A2(_1459_),
    .A3(_1477_),
    .B1(_1479_),
    .X(_0319_));
 sky130_fd_sc_hd__or2b_1 _4070_ (.A(_1457_),
    .B_N(_1456_),
    .X(_1480_));
 sky130_fd_sc_hd__nand2_1 _4071_ (.A(_1292_),
    .B(_1453_),
    .Y(_1481_));
 sky130_fd_sc_hd__xnor2_1 _4072_ (.A(_1480_),
    .B(_1481_),
    .Y(_1482_));
 sky130_fd_sc_hd__mux2_1 _4073_ (.A0(net563),
    .A1(_1482_),
    .S(_1468_),
    .X(_1483_));
 sky130_fd_sc_hd__or4_4 _4074_ (.A(net265),
    .B(net262),
    .C(net261),
    .D(_0870_),
    .X(_1484_));
 sky130_fd_sc_hd__nand2_4 _4075_ (.A(_1484_),
    .B(_0999_),
    .Y(_1485_));
 sky130_fd_sc_hd__mux2_1 _4076_ (.A0(net324),
    .A1(_1483_),
    .S(_1485_),
    .X(_1486_));
 sky130_fd_sc_hd__clkbuf_1 _4077_ (.A(_1486_),
    .X(_0318_));
 sky130_fd_sc_hd__buf_2 _4078_ (.A(_0999_),
    .X(_1487_));
 sky130_fd_sc_hd__clkbuf_2 _4079_ (.A(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__buf_2 _4080_ (.A(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__mux2_1 _4081_ (.A0(net325),
    .A1(net541),
    .S(_0893_),
    .X(_1490_));
 sky130_fd_sc_hd__buf_2 _4082_ (.A(_1468_),
    .X(_1491_));
 sky130_fd_sc_hd__nand3_1 _4083_ (.A(_1452_),
    .B(_1443_),
    .C(_1451_),
    .Y(_1492_));
 sky130_fd_sc_hd__and3_1 _4084_ (.A(_1491_),
    .B(_1453_),
    .C(_1492_),
    .X(_1493_));
 sky130_fd_sc_hd__a21o_1 _4085_ (.A1(_1489_),
    .A2(_1490_),
    .B1(_1493_),
    .X(_0317_));
 sky130_fd_sc_hd__inv_2 _4086_ (.A(net569),
    .Y(_1494_));
 sky130_fd_sc_hd__a21oi_1 _4087_ (.A1(_1414_),
    .A2(_1426_),
    .B1(_1432_),
    .Y(_1495_));
 sky130_fd_sc_hd__o21ai_1 _4088_ (.A1(_1495_),
    .A2(_1447_),
    .B1(_1445_),
    .Y(_1496_));
 sky130_fd_sc_hd__nor2_1 _4089_ (.A(_1441_),
    .B(_1496_),
    .Y(_1497_));
 sky130_fd_sc_hd__o21ai_1 _4090_ (.A1(_1448_),
    .A2(_1497_),
    .B1(_1439_),
    .Y(_1498_));
 sky130_fd_sc_hd__o31a_1 _4091_ (.A1(_1439_),
    .A2(_1448_),
    .A3(_1497_),
    .B1(_1468_),
    .X(_1499_));
 sky130_fd_sc_hd__a221o_1 _4092_ (.A1(_1494_),
    .A2(_1488_),
    .B1(_1498_),
    .B2(_1499_),
    .C1(_1473_),
    .X(_1500_));
 sky130_fd_sc_hd__a21bo_1 _4093_ (.A1(net326),
    .A2(_1474_),
    .B1_N(_1500_),
    .X(_0316_));
 sky130_fd_sc_hd__clkbuf_2 _4094_ (.A(_1473_),
    .X(_1501_));
 sky130_fd_sc_hd__or2_1 _4095_ (.A(_1487_),
    .B(_1497_),
    .X(_1502_));
 sky130_fd_sc_hd__a21oi_1 _4096_ (.A1(_1441_),
    .A2(_1496_),
    .B1(_1502_),
    .Y(_1503_));
 sky130_fd_sc_hd__a221o_1 _4097_ (.A1(net457),
    .A2(_0894_),
    .B1(_1501_),
    .B2(net329),
    .C1(_1503_),
    .X(_0315_));
 sky130_fd_sc_hd__o21bai_1 _4098_ (.A1(_1430_),
    .A2(_1495_),
    .B1_N(_1436_),
    .Y(_1504_));
 sky130_fd_sc_hd__or3b_1 _4099_ (.A(_1430_),
    .B(_1495_),
    .C_N(_1436_),
    .X(_1505_));
 sky130_fd_sc_hd__a22o_1 _4100_ (.A1(net498),
    .A2(_0880_),
    .B1(_1473_),
    .B2(net331),
    .X(_1506_));
 sky130_fd_sc_hd__a31o_1 _4101_ (.A1(_1475_),
    .A2(_1504_),
    .A3(_1505_),
    .B1(_1506_),
    .X(_0314_));
 sky130_fd_sc_hd__and3_1 _4102_ (.A(_1414_),
    .B(_1426_),
    .C(_1432_),
    .X(_1507_));
 sky130_fd_sc_hd__nor2_1 _4103_ (.A(_1495_),
    .B(_1507_),
    .Y(_1508_));
 sky130_fd_sc_hd__a22o_1 _4104_ (.A1(net515),
    .A2(_0889_),
    .B1(_1478_),
    .B2(net333),
    .X(_1509_));
 sky130_fd_sc_hd__a21o_1 _4105_ (.A1(_1475_),
    .A2(_1508_),
    .B1(_1509_),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_2 _4106_ (.A(_1485_),
    .X(_1510_));
 sky130_fd_sc_hd__a21oi_1 _4107_ (.A1(_1294_),
    .A2(_1374_),
    .B1(_1393_),
    .Y(_1511_));
 sky130_fd_sc_hd__a221o_1 _4108_ (.A1(net341),
    .A2(_1376_),
    .B1(_1415_),
    .B2(_1416_),
    .C1(_1417_),
    .X(_1512_));
 sky130_fd_sc_hd__o21a_1 _4109_ (.A1(_1511_),
    .A2(_1512_),
    .B1(_1406_),
    .X(_1513_));
 sky130_fd_sc_hd__or3_1 _4110_ (.A(_1404_),
    .B(_1411_),
    .C(_1513_),
    .X(_1514_));
 sky130_fd_sc_hd__a31o_1 _4111_ (.A1(_1399_),
    .A2(_1419_),
    .A3(_1514_),
    .B1(_1423_),
    .X(_1515_));
 sky130_fd_sc_hd__xnor2_1 _4112_ (.A(_1396_),
    .B(_1515_),
    .Y(_1516_));
 sky130_fd_sc_hd__nor2_1 _4113_ (.A(net545),
    .B(_1491_),
    .Y(_1517_));
 sky130_fd_sc_hd__a211o_1 _4114_ (.A1(_1491_),
    .A2(_1516_),
    .B1(_1517_),
    .C1(_1478_),
    .X(_1518_));
 sky130_fd_sc_hd__o21ai_1 _4115_ (.A1(_1421_),
    .A2(_1510_),
    .B1(_1518_),
    .Y(_0312_));
 sky130_fd_sc_hd__a21oi_1 _4116_ (.A1(_1419_),
    .A2(_1514_),
    .B1(_1399_),
    .Y(_1519_));
 sky130_fd_sc_hd__a31o_1 _4117_ (.A1(_1399_),
    .A2(_1419_),
    .A3(_1514_),
    .B1(_1487_),
    .X(_1520_));
 sky130_fd_sc_hd__nor2_1 _4118_ (.A(_1519_),
    .B(_1520_),
    .Y(_1521_));
 sky130_fd_sc_hd__a221o_1 _4119_ (.A1(net467),
    .A2(_0949_),
    .B1(_1474_),
    .B2(net337),
    .C1(_1521_),
    .X(_0311_));
 sky130_fd_sc_hd__nor2_1 _4120_ (.A(_1404_),
    .B(_1513_),
    .Y(_1522_));
 sky130_fd_sc_hd__xnor2_1 _4121_ (.A(_1412_),
    .B(_1522_),
    .Y(_1523_));
 sky130_fd_sc_hd__mux2_1 _4122_ (.A0(net559),
    .A1(_1523_),
    .S(_1153_),
    .X(_1524_));
 sky130_fd_sc_hd__mux2_1 _4123_ (.A0(net338),
    .A1(_1524_),
    .S(_1485_),
    .X(_1525_));
 sky130_fd_sc_hd__clkbuf_1 _4124_ (.A(_1525_),
    .X(_0310_));
 sky130_fd_sc_hd__nor2_1 _4125_ (.A(_1487_),
    .B(_1513_),
    .Y(_1526_));
 sky130_fd_sc_hd__o31a_1 _4126_ (.A1(_1406_),
    .A2(_1511_),
    .A3(_1512_),
    .B1(_1526_),
    .X(_1527_));
 sky130_fd_sc_hd__a221o_1 _4127_ (.A1(net459),
    .A2(_0902_),
    .B1(_1474_),
    .B2(net340),
    .C1(_1527_),
    .X(_0309_));
 sky130_fd_sc_hd__a21o_1 _4128_ (.A1(net539),
    .A2(_0949_),
    .B1(_1469_),
    .X(_1528_));
 sky130_fd_sc_hd__or2_1 _4129_ (.A(_1380_),
    .B(_1381_),
    .X(_1529_));
 sky130_fd_sc_hd__a21oi_2 _4130_ (.A1(_1294_),
    .A2(_1374_),
    .B1(_1392_),
    .Y(_1530_));
 sky130_fd_sc_hd__o21bai_1 _4131_ (.A1(_1416_),
    .A2(_1530_),
    .B1_N(_1385_),
    .Y(_1531_));
 sky130_fd_sc_hd__o21ba_1 _4132_ (.A1(_1529_),
    .A2(_1531_),
    .B1_N(_1380_),
    .X(_1532_));
 sky130_fd_sc_hd__xnor2_1 _4133_ (.A(_1377_),
    .B(_1532_),
    .Y(_1533_));
 sky130_fd_sc_hd__nand2_1 _4134_ (.A(_1469_),
    .B(_1533_),
    .Y(_1534_));
 sky130_fd_sc_hd__a22o_1 _4135_ (.A1(net343),
    .A2(_1474_),
    .B1(_1528_),
    .B2(_1534_),
    .X(_0308_));
 sky130_fd_sc_hd__o21ai_1 _4136_ (.A1(_1529_),
    .A2(_1531_),
    .B1(_1491_),
    .Y(_1535_));
 sky130_fd_sc_hd__a21oi_1 _4137_ (.A1(_1529_),
    .A2(_1531_),
    .B1(_1535_),
    .Y(_1536_));
 sky130_fd_sc_hd__a221o_1 _4138_ (.A1(net475),
    .A2(_0949_),
    .B1(_1478_),
    .B2(net345),
    .C1(_1536_),
    .X(_0307_));
 sky130_fd_sc_hd__nor2_1 _4139_ (.A(_1385_),
    .B(_1387_),
    .Y(_1537_));
 sky130_fd_sc_hd__o21ai_1 _4140_ (.A1(_1391_),
    .A2(_1530_),
    .B1(_1537_),
    .Y(_1538_));
 sky130_fd_sc_hd__o311a_1 _4141_ (.A1(_1391_),
    .A2(_1530_),
    .A3(_1537_),
    .B1(_1538_),
    .C1(_1491_),
    .X(_1539_));
 sky130_fd_sc_hd__a221o_1 _4142_ (.A1(net453),
    .A2(_0902_),
    .B1(_1501_),
    .B2(net347),
    .C1(_1539_),
    .X(_0306_));
 sky130_fd_sc_hd__and3_1 _4143_ (.A(_1294_),
    .B(_1374_),
    .C(_1392_),
    .X(_1540_));
 sky130_fd_sc_hd__nor3_1 _4144_ (.A(_1488_),
    .B(_1530_),
    .C(_1540_),
    .Y(_1541_));
 sky130_fd_sc_hd__a221o_1 _4145_ (.A1(net461),
    .A2(_0949_),
    .B1(_1478_),
    .B2(net349),
    .C1(_1541_),
    .X(_0305_));
 sky130_fd_sc_hd__clkbuf_2 _4146_ (.A(_1484_),
    .X(_1542_));
 sky130_fd_sc_hd__or3_1 _4147_ (.A(_1373_),
    .B(_1297_),
    .C(_1371_),
    .X(_1543_));
 sky130_fd_sc_hd__a21o_1 _4148_ (.A1(_1374_),
    .A2(_1543_),
    .B1(_1488_),
    .X(_1544_));
 sky130_fd_sc_hd__o221a_1 _4149_ (.A1(net479),
    .A2(_1542_),
    .B1(_1510_),
    .B2(net351),
    .C1(_1544_),
    .X(_0304_));
 sky130_fd_sc_hd__a311oi_1 _4150_ (.A1(_1370_),
    .A2(_1305_),
    .A3(_1367_),
    .B1(_1371_),
    .C1(_1488_),
    .Y(_1545_));
 sky130_fd_sc_hd__a221o_1 _4151_ (.A1(net477),
    .A2(_0894_),
    .B1(_1501_),
    .B2(net353),
    .C1(_1545_),
    .X(_0303_));
 sky130_fd_sc_hd__o31ai_1 _4152_ (.A1(_1307_),
    .A2(_1310_),
    .A3(_1365_),
    .B1(_1303_),
    .Y(_1546_));
 sky130_fd_sc_hd__xnor2_1 _4153_ (.A(_1546_),
    .B(_1366_),
    .Y(_1547_));
 sky130_fd_sc_hd__mux2_1 _4154_ (.A0(net567),
    .A1(_1547_),
    .S(_1468_),
    .X(_1548_));
 sky130_fd_sc_hd__mux2_1 _4155_ (.A0(net355),
    .A1(_1548_),
    .S(_1485_),
    .X(_1549_));
 sky130_fd_sc_hd__clkbuf_1 _4156_ (.A(_1549_),
    .X(_0302_));
 sky130_fd_sc_hd__nor2_1 _4157_ (.A(_1310_),
    .B(_1365_),
    .Y(_1550_));
 sky130_fd_sc_hd__xnor2_1 _4158_ (.A(_1307_),
    .B(_1550_),
    .Y(_1551_));
 sky130_fd_sc_hd__or2_1 _4159_ (.A(net543),
    .B(_1542_),
    .X(_1552_));
 sky130_fd_sc_hd__o221a_1 _4160_ (.A1(net357),
    .A2(_1510_),
    .B1(_1551_),
    .B2(_1489_),
    .C1(_1552_),
    .X(_0301_));
 sky130_fd_sc_hd__o31a_1 _4161_ (.A1(_1313_),
    .A2(_1357_),
    .A3(_1363_),
    .B1(_1360_),
    .X(_1553_));
 sky130_fd_sc_hd__and2b_1 _4162_ (.A_N(_1310_),
    .B(_1364_),
    .X(_1554_));
 sky130_fd_sc_hd__xnor2_1 _4163_ (.A(_1553_),
    .B(_1554_),
    .Y(_1555_));
 sky130_fd_sc_hd__mux2_1 _4164_ (.A0(net561),
    .A1(_1555_),
    .S(_1153_),
    .X(_1556_));
 sky130_fd_sc_hd__mux2_1 _4165_ (.A0(net358),
    .A1(_1556_),
    .S(_1485_),
    .X(_1557_));
 sky130_fd_sc_hd__clkbuf_1 _4166_ (.A(_1557_),
    .X(_0300_));
 sky130_fd_sc_hd__nor2_1 _4167_ (.A(_1313_),
    .B(_1357_),
    .Y(_1558_));
 sky130_fd_sc_hd__xnor2_1 _4168_ (.A(_1558_),
    .B(_1363_),
    .Y(_1559_));
 sky130_fd_sc_hd__or2_1 _4169_ (.A(net549),
    .B(_1542_),
    .X(_1560_));
 sky130_fd_sc_hd__o221a_1 _4170_ (.A1(net361),
    .A2(_1510_),
    .B1(_1559_),
    .B2(_1489_),
    .C1(_1560_),
    .X(_0299_));
 sky130_fd_sc_hd__or2_1 _4171_ (.A(_1319_),
    .B(_1354_),
    .X(_1561_));
 sky130_fd_sc_hd__nand2_1 _4172_ (.A(_1316_),
    .B(_1561_),
    .Y(_1562_));
 sky130_fd_sc_hd__o21ai_1 _4173_ (.A1(_1313_),
    .A2(_1355_),
    .B1(_1562_),
    .Y(_1563_));
 sky130_fd_sc_hd__o31a_1 _4174_ (.A1(_1313_),
    .A2(_1355_),
    .A3(_1562_),
    .B1(_1468_),
    .X(_1564_));
 sky130_fd_sc_hd__nand2_1 _4175_ (.A(_1563_),
    .B(_1564_),
    .Y(_1565_));
 sky130_fd_sc_hd__a21o_1 _4176_ (.A1(net537),
    .A2(_0889_),
    .B1(_1469_),
    .X(_1566_));
 sky130_fd_sc_hd__a22o_1 _4177_ (.A1(net362),
    .A2(_1474_),
    .B1(_1565_),
    .B2(_1566_),
    .X(_0298_));
 sky130_fd_sc_hd__nand2_1 _4178_ (.A(_1319_),
    .B(_1354_),
    .Y(_1567_));
 sky130_fd_sc_hd__a22o_1 _4179_ (.A1(net504),
    .A2(_0874_),
    .B1(_1478_),
    .B2(net364),
    .X(_1568_));
 sky130_fd_sc_hd__a31o_1 _4180_ (.A1(_1475_),
    .A2(_1561_),
    .A3(_1567_),
    .B1(_1568_),
    .X(_0297_));
 sky130_fd_sc_hd__and2b_1 _4181_ (.A_N(_1353_),
    .B(_1322_),
    .X(_1569_));
 sky130_fd_sc_hd__a21oi_1 _4182_ (.A1(_1569_),
    .A2(_1352_),
    .B1(_1487_),
    .Y(_1570_));
 sky130_fd_sc_hd__o21a_1 _4183_ (.A1(_1569_),
    .A2(_1352_),
    .B1(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__a221o_1 _4184_ (.A1(net449),
    .A2(_0894_),
    .B1(_1501_),
    .B2(net366),
    .C1(_1571_),
    .X(_0296_));
 sky130_fd_sc_hd__nand2_1 _4185_ (.A(_1325_),
    .B(_1350_),
    .Y(_1572_));
 sky130_fd_sc_hd__or2_1 _4186_ (.A(_1325_),
    .B(_1350_),
    .X(_1573_));
 sky130_fd_sc_hd__a22o_1 _4187_ (.A1(net494),
    .A2(_0880_),
    .B1(_1473_),
    .B2(net368),
    .X(_1574_));
 sky130_fd_sc_hd__a31o_1 _4188_ (.A1(_1475_),
    .A2(_1572_),
    .A3(_1573_),
    .B1(_1574_),
    .X(_0295_));
 sky130_fd_sc_hd__xor2_1 _4189_ (.A(_1330_),
    .B(_1348_),
    .X(_1575_));
 sky130_fd_sc_hd__or2_1 _4190_ (.A(net553),
    .B(_1484_),
    .X(_1576_));
 sky130_fd_sc_hd__o221a_1 _4191_ (.A1(net371),
    .A2(_1510_),
    .B1(_1575_),
    .B2(_1489_),
    .C1(_1576_),
    .X(_0294_));
 sky130_fd_sc_hd__xor2_1 _4192_ (.A(_1344_),
    .B(_1346_),
    .X(_1577_));
 sky130_fd_sc_hd__or2_1 _4193_ (.A(net547),
    .B(_1542_),
    .X(_1578_));
 sky130_fd_sc_hd__o221a_1 _4194_ (.A1(net372),
    .A2(_1510_),
    .B1(_1577_),
    .B2(_1489_),
    .C1(_1578_),
    .X(_0293_));
 sky130_fd_sc_hd__nand2_1 _4195_ (.A(_1332_),
    .B(_1342_),
    .Y(_1579_));
 sky130_fd_sc_hd__or2_1 _4196_ (.A(_1332_),
    .B(_1342_),
    .X(_1580_));
 sky130_fd_sc_hd__and3_1 _4197_ (.A(_1491_),
    .B(_1579_),
    .C(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__a221o_1 _4198_ (.A1(net455),
    .A2(_0894_),
    .B1(_1501_),
    .B2(net373),
    .C1(_1581_),
    .X(_0292_));
 sky130_fd_sc_hd__and2b_1 _4199_ (.A_N(_1341_),
    .B(_1340_),
    .X(_1582_));
 sky130_fd_sc_hd__xnor2_1 _4200_ (.A(_1337_),
    .B(_1582_),
    .Y(_1583_));
 sky130_fd_sc_hd__nor2_1 _4201_ (.A(_1488_),
    .B(_1583_),
    .Y(_1584_));
 sky130_fd_sc_hd__a221o_1 _4202_ (.A1(net451),
    .A2(_0894_),
    .B1(_1501_),
    .B2(net374),
    .C1(_1584_),
    .X(_0291_));
 sky130_fd_sc_hd__nand2_1 _4203_ (.A(net376),
    .B(_1198_),
    .Y(_1585_));
 sky130_fd_sc_hd__or2b_1 _4204_ (.A(_1336_),
    .B_N(_1335_),
    .X(_1586_));
 sky130_fd_sc_hd__or2_1 _4205_ (.A(_1585_),
    .B(_1586_),
    .X(_1587_));
 sky130_fd_sc_hd__nand2_1 _4206_ (.A(_1585_),
    .B(_1586_),
    .Y(_1588_));
 sky130_fd_sc_hd__a22o_1 _4207_ (.A1(net517),
    .A2(_0874_),
    .B1(_1473_),
    .B2(net375),
    .X(_1589_));
 sky130_fd_sc_hd__a31o_1 _4208_ (.A1(_1475_),
    .A2(_1587_),
    .A3(_1588_),
    .B1(_1589_),
    .X(_0290_));
 sky130_fd_sc_hd__o21a_1 _4209_ (.A1(_1487_),
    .A2(_1198_),
    .B1(_1485_),
    .X(_1590_));
 sky130_fd_sc_hd__o22a_1 _4210_ (.A1(net555),
    .A2(_1542_),
    .B1(_1590_),
    .B2(net376),
    .X(_1591_));
 sky130_fd_sc_hd__o21a_1 _4211_ (.A1(_1489_),
    .A2(_1585_),
    .B1(net556),
    .X(_0289_));
 sky130_fd_sc_hd__or4_1 _4212_ (.A(\state[4] ),
    .B(net264),
    .C(_0867_),
    .D(_0769_),
    .X(_1592_));
 sky130_fd_sc_hd__nor2_2 _4213_ (.A(\state[0] ),
    .B(_1592_),
    .Y(_1593_));
 sky130_fd_sc_hd__nor2_1 _4214_ (.A(_0997_),
    .B(_0870_),
    .Y(_1594_));
 sky130_fd_sc_hd__and3_1 _4215_ (.A(net262),
    .B(_0769_),
    .C(_1594_),
    .X(_1595_));
 sky130_fd_sc_hd__nor2_1 _4216_ (.A(_1593_),
    .B(_1595_),
    .Y(_1596_));
 sky130_fd_sc_hd__nand2_1 _4217_ (.A(_1484_),
    .B(_1596_),
    .Y(_1597_));
 sky130_fd_sc_hd__buf_2 _4218_ (.A(_1597_),
    .X(_1598_));
 sky130_fd_sc_hd__and4bb_1 _4219_ (.A_N(\state[4] ),
    .B_N(net265),
    .C(net262),
    .D(net261),
    .X(_1599_));
 sky130_fd_sc_hd__inv_2 _4220_ (.A(net398),
    .Y(_1600_));
 sky130_fd_sc_hd__a21oi_1 _4221_ (.A1(_0868_),
    .A2(_1599_),
    .B1(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__clkbuf_2 _4222_ (.A(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__clkbuf_2 _4223_ (.A(_1602_),
    .X(_1603_));
 sky130_fd_sc_hd__clkbuf_2 _4224_ (.A(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4225_ (.A(_1604_),
    .X(_1605_));
 sky130_fd_sc_hd__or2_1 _4226_ (.A(\sum[30] ),
    .B(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__or2_1 _4227_ (.A(\sum[29] ),
    .B(_1605_),
    .X(_1607_));
 sky130_fd_sc_hd__and3_1 _4228_ (.A(net398),
    .B(_0868_),
    .C(_1599_),
    .X(_1608_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4229_ (.A(_1608_),
    .X(_1609_));
 sky130_fd_sc_hd__buf_1 _4230_ (.A(_1609_),
    .X(_1610_));
 sky130_fd_sc_hd__buf_1 _4231_ (.A(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__buf_1 _4232_ (.A(_1611_),
    .X(_1612_));
 sky130_fd_sc_hd__buf_2 _4233_ (.A(_1612_),
    .X(_1613_));
 sky130_fd_sc_hd__clkbuf_2 _4234_ (.A(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__xor2_1 _4235_ (.A(\sum[27] ),
    .B(_1614_),
    .X(_1615_));
 sky130_fd_sc_hd__and2_1 _4236_ (.A(\sum[17] ),
    .B(_1612_),
    .X(_1616_));
 sky130_fd_sc_hd__and2_1 _4237_ (.A(\sum[16] ),
    .B(_1612_),
    .X(_1617_));
 sky130_fd_sc_hd__and2_1 _4238_ (.A(\sum[14] ),
    .B(_1610_),
    .X(_1618_));
 sky130_fd_sc_hd__o21a_1 _4239_ (.A1(_1603_),
    .A2(_1618_),
    .B1(\sum[15] ),
    .X(_1619_));
 sky130_fd_sc_hd__and2_1 _4240_ (.A(net380),
    .B(_1610_),
    .X(_1620_));
 sky130_fd_sc_hd__and2_1 _4241_ (.A(\sum[10] ),
    .B(_1602_),
    .X(_1621_));
 sky130_fd_sc_hd__nor2_1 _4242_ (.A(\sum[10] ),
    .B(_1603_),
    .Y(_1622_));
 sky130_fd_sc_hd__or2_1 _4243_ (.A(_1621_),
    .B(_1622_),
    .X(_1623_));
 sky130_fd_sc_hd__or2_1 _4244_ (.A(net382),
    .B(_1603_),
    .X(_1624_));
 sky130_fd_sc_hd__or2_1 _4245_ (.A(\sum[7] ),
    .B(_1609_),
    .X(_1625_));
 sky130_fd_sc_hd__nor2_1 _4246_ (.A(net383),
    .B(_1602_),
    .Y(_1626_));
 sky130_fd_sc_hd__nor2_1 _4247_ (.A(\sum[5] ),
    .B(_1609_),
    .Y(_1627_));
 sky130_fd_sc_hd__or2_1 _4248_ (.A(\sum[3] ),
    .B(_1608_),
    .X(_1628_));
 sky130_fd_sc_hd__or2_1 _4249_ (.A(net384),
    .B(_1601_),
    .X(_1629_));
 sky130_fd_sc_hd__and2_1 _4250_ (.A(net384),
    .B(_1601_),
    .X(_1630_));
 sky130_fd_sc_hd__a31o_1 _4251_ (.A1(\sum[0] ),
    .A2(net398),
    .A3(_1629_),
    .B1(_1630_),
    .X(_1631_));
 sky130_fd_sc_hd__or2_1 _4252_ (.A(\sum[2] ),
    .B(_1601_),
    .X(_1632_));
 sky130_fd_sc_hd__and2_1 _4253_ (.A(\sum[2] ),
    .B(_1602_),
    .X(_1633_));
 sky130_fd_sc_hd__a21o_1 _4254_ (.A1(_1631_),
    .A2(_1632_),
    .B1(_1633_),
    .X(_1634_));
 sky130_fd_sc_hd__nand2_1 _4255_ (.A(\sum[3] ),
    .B(_1608_),
    .Y(_1635_));
 sky130_fd_sc_hd__a21bo_1 _4256_ (.A1(_1628_),
    .A2(_1634_),
    .B1_N(_1635_),
    .X(_1636_));
 sky130_fd_sc_hd__and2_1 _4257_ (.A(\sum[4] ),
    .B(_1608_),
    .X(_1637_));
 sky130_fd_sc_hd__nor2_1 _4258_ (.A(\sum[4] ),
    .B(_1608_),
    .Y(_1638_));
 sky130_fd_sc_hd__nor2_1 _4259_ (.A(_1637_),
    .B(_1638_),
    .Y(_1639_));
 sky130_fd_sc_hd__and2_1 _4260_ (.A(\sum[5] ),
    .B(_1608_),
    .X(_1640_));
 sky130_fd_sc_hd__a211oi_2 _4261_ (.A1(_1636_),
    .A2(_1639_),
    .B1(_1640_),
    .C1(_1637_),
    .Y(_1641_));
 sky130_fd_sc_hd__nand2_1 _4262_ (.A(\sum[6] ),
    .B(_1602_),
    .Y(_1642_));
 sky130_fd_sc_hd__o31ai_2 _4263_ (.A1(_1626_),
    .A2(_1627_),
    .A3(_1641_),
    .B1(_1642_),
    .Y(_1643_));
 sky130_fd_sc_hd__nand2_1 _4264_ (.A(\sum[7] ),
    .B(_1609_),
    .Y(_1644_));
 sky130_fd_sc_hd__a21bo_1 _4265_ (.A1(_1625_),
    .A2(_1643_),
    .B1_N(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__or2_1 _4266_ (.A(\sum[8] ),
    .B(_1609_),
    .X(_1646_));
 sky130_fd_sc_hd__and2_1 _4267_ (.A(net382),
    .B(_1602_),
    .X(_1647_));
 sky130_fd_sc_hd__and2_1 _4268_ (.A(\sum[8] ),
    .B(_1609_),
    .X(_1648_));
 sky130_fd_sc_hd__a211o_1 _4269_ (.A1(_1645_),
    .A2(_1646_),
    .B1(_1647_),
    .C1(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__and3b_1 _4270_ (.A_N(_1623_),
    .B(_1624_),
    .C(_1649_),
    .X(_1650_));
 sky130_fd_sc_hd__nand2_1 _4271_ (.A(net379),
    .B(_1610_),
    .Y(_1651_));
 sky130_fd_sc_hd__or2_1 _4272_ (.A(net379),
    .B(_1610_),
    .X(_1652_));
 sky130_fd_sc_hd__nand2_1 _4273_ (.A(_1651_),
    .B(_1652_),
    .Y(_1653_));
 sky130_fd_sc_hd__inv_2 _4274_ (.A(_1653_),
    .Y(_1654_));
 sky130_fd_sc_hd__or2_1 _4275_ (.A(net380),
    .B(_1611_),
    .X(_1655_));
 sky130_fd_sc_hd__o311a_1 _4276_ (.A1(_1620_),
    .A2(_1621_),
    .A3(_1650_),
    .B1(_1654_),
    .C1(_1655_),
    .X(_1656_));
 sky130_fd_sc_hd__nand2_1 _4277_ (.A(\sum[13] ),
    .B(_1611_),
    .Y(_1657_));
 sky130_fd_sc_hd__nand2_1 _4278_ (.A(_1657_),
    .B(_1651_),
    .Y(_1658_));
 sky130_fd_sc_hd__or2_1 _4279_ (.A(\sum[15] ),
    .B(_1603_),
    .X(_1659_));
 sky130_fd_sc_hd__nor2_1 _4280_ (.A(\sum[14] ),
    .B(_1610_),
    .Y(_1660_));
 sky130_fd_sc_hd__or2_1 _4281_ (.A(_1618_),
    .B(_1660_),
    .X(_1661_));
 sky130_fd_sc_hd__inv_2 _4282_ (.A(_1661_),
    .Y(_1662_));
 sky130_fd_sc_hd__or2_1 _4283_ (.A(\sum[13] ),
    .B(_1611_),
    .X(_1663_));
 sky130_fd_sc_hd__o2111a_1 _4284_ (.A1(_1656_),
    .A2(_1658_),
    .B1(_1659_),
    .C1(_1662_),
    .D1(_1663_),
    .X(_1664_));
 sky130_fd_sc_hd__or2_1 _4285_ (.A(\sum[16] ),
    .B(_1612_),
    .X(_1665_));
 sky130_fd_sc_hd__nand2_1 _4286_ (.A(\sum[16] ),
    .B(_1612_),
    .Y(_1666_));
 sky130_fd_sc_hd__o211a_1 _4287_ (.A1(_1619_),
    .A2(_1664_),
    .B1(_1665_),
    .C1(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__or2_1 _4288_ (.A(\sum[17] ),
    .B(_1612_),
    .X(_1668_));
 sky130_fd_sc_hd__and2_1 _4289_ (.A(\sum[18] ),
    .B(_1611_),
    .X(_1669_));
 sky130_fd_sc_hd__nor2_1 _4290_ (.A(\sum[18] ),
    .B(_1611_),
    .Y(_1670_));
 sky130_fd_sc_hd__or2_1 _4291_ (.A(_1669_),
    .B(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__inv_2 _4292_ (.A(_1671_),
    .Y(_1672_));
 sky130_fd_sc_hd__o311a_1 _4293_ (.A1(_1616_),
    .A2(_1617_),
    .A3(_1667_),
    .B1(_1668_),
    .C1(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__or2_1 _4294_ (.A(net378),
    .B(_1604_),
    .X(_1674_));
 sky130_fd_sc_hd__o21a_1 _4295_ (.A1(_1604_),
    .A2(_1669_),
    .B1(net378),
    .X(_1675_));
 sky130_fd_sc_hd__a21oi_1 _4296_ (.A1(_1673_),
    .A2(_1674_),
    .B1(_1675_),
    .Y(_1676_));
 sky130_fd_sc_hd__xnor2_1 _4297_ (.A(\sum[20] ),
    .B(_1613_),
    .Y(_1677_));
 sky130_fd_sc_hd__and2_1 _4298_ (.A(\sum[22] ),
    .B(_1603_),
    .X(_1678_));
 sky130_fd_sc_hd__nor2_1 _4299_ (.A(\sum[22] ),
    .B(_1604_),
    .Y(_1679_));
 sky130_fd_sc_hd__or2_1 _4300_ (.A(_1678_),
    .B(_1679_),
    .X(_1680_));
 sky130_fd_sc_hd__xnor2_1 _4301_ (.A(\sum[23] ),
    .B(_1604_),
    .Y(_1681_));
 sky130_fd_sc_hd__nor2_1 _4302_ (.A(_1680_),
    .B(_1681_),
    .Y(_1682_));
 sky130_fd_sc_hd__xnor2_1 _4303_ (.A(\sum[21] ),
    .B(_1613_),
    .Y(_1683_));
 sky130_fd_sc_hd__inv_2 _4304_ (.A(_1683_),
    .Y(_1684_));
 sky130_fd_sc_hd__and4bb_1 _4305_ (.A_N(_1676_),
    .B_N(_1677_),
    .C(_1682_),
    .D(_1684_),
    .X(_1685_));
 sky130_fd_sc_hd__o21a_1 _4306_ (.A1(\sum[21] ),
    .A2(\sum[20] ),
    .B1(_1613_),
    .X(_1686_));
 sky130_fd_sc_hd__o21a_1 _4307_ (.A1(\sum[23] ),
    .A2(\sum[22] ),
    .B1(_1604_),
    .X(_1687_));
 sky130_fd_sc_hd__a21o_1 _4308_ (.A1(_1682_),
    .A2(_1686_),
    .B1(_1687_),
    .X(_1688_));
 sky130_fd_sc_hd__xor2_1 _4309_ (.A(\sum[24] ),
    .B(_1605_),
    .X(_1689_));
 sky130_fd_sc_hd__o21ai_1 _4310_ (.A1(_1685_),
    .A2(_1688_),
    .B1(_1689_),
    .Y(_1690_));
 sky130_fd_sc_hd__xnor2_1 _4311_ (.A(\sum[25] ),
    .B(_1613_),
    .Y(_1691_));
 sky130_fd_sc_hd__or2_1 _4312_ (.A(_1690_),
    .B(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__o211ai_1 _4313_ (.A1(\sum[24] ),
    .A2(_1593_),
    .B1(net399),
    .C1(\sum[25] ),
    .Y(_1693_));
 sky130_fd_sc_hd__xnor2_1 _4314_ (.A(\sum[26] ),
    .B(_1613_),
    .Y(_1694_));
 sky130_fd_sc_hd__a21oi_1 _4315_ (.A1(_1692_),
    .A2(_1693_),
    .B1(_1694_),
    .Y(_1695_));
 sky130_fd_sc_hd__o21a_1 _4316_ (.A1(\sum[27] ),
    .A2(\sum[26] ),
    .B1(_1614_),
    .X(_1696_));
 sky130_fd_sc_hd__a21oi_1 _4317_ (.A1(_1615_),
    .A2(_1695_),
    .B1(_1696_),
    .Y(_1697_));
 sky130_fd_sc_hd__xnor2_1 _4318_ (.A(\sum[28] ),
    .B(_1614_),
    .Y(_1698_));
 sky130_fd_sc_hd__a2bb2o_1 _4319_ (.A1_N(_1697_),
    .A2_N(_1698_),
    .B1(\sum[28] ),
    .B2(_1614_),
    .X(_1699_));
 sky130_fd_sc_hd__nand2_1 _4320_ (.A(\sum[29] ),
    .B(_1605_),
    .Y(_1700_));
 sky130_fd_sc_hd__a21bo_1 _4321_ (.A1(_1607_),
    .A2(_1699_),
    .B1_N(_1700_),
    .X(_1701_));
 sky130_fd_sc_hd__and2_1 _4322_ (.A(\sum[30] ),
    .B(_1605_),
    .X(_1702_));
 sky130_fd_sc_hd__a21o_1 _4323_ (.A1(_1606_),
    .A2(_1701_),
    .B1(_1702_),
    .X(_1703_));
 sky130_fd_sc_hd__buf_2 _4324_ (.A(_1614_),
    .X(_1704_));
 sky130_fd_sc_hd__xnor2_1 _4325_ (.A(\sum[31] ),
    .B(_1704_),
    .Y(_1705_));
 sky130_fd_sc_hd__xnor2_1 _4326_ (.A(_1703_),
    .B(_1705_),
    .Y(_1706_));
 sky130_fd_sc_hd__buf_2 _4327_ (.A(_1596_),
    .X(_1707_));
 sky130_fd_sc_hd__buf_2 _4328_ (.A(_1707_),
    .X(_1708_));
 sky130_fd_sc_hd__o22a_1 _4329_ (.A1(\sum[31] ),
    .A2(_1598_),
    .B1(_1706_),
    .B2(_1708_),
    .X(_0288_));
 sky130_fd_sc_hd__or2b_1 _4330_ (.A(_1702_),
    .B_N(_1606_),
    .X(_1709_));
 sky130_fd_sc_hd__xnor2_1 _4331_ (.A(_1709_),
    .B(_1701_),
    .Y(_1710_));
 sky130_fd_sc_hd__buf_2 _4332_ (.A(_1707_),
    .X(_1711_));
 sky130_fd_sc_hd__o22a_1 _4333_ (.A1(\sum[30] ),
    .A2(_1598_),
    .B1(_1710_),
    .B2(_1711_),
    .X(_0287_));
 sky130_fd_sc_hd__or2_1 _4334_ (.A(_1593_),
    .B(_1595_),
    .X(_1712_));
 sky130_fd_sc_hd__nor2_2 _4335_ (.A(_0893_),
    .B(_1712_),
    .Y(_1713_));
 sky130_fd_sc_hd__buf_2 _4336_ (.A(_1713_),
    .X(_1714_));
 sky130_fd_sc_hd__nand2_1 _4337_ (.A(_1607_),
    .B(_1700_),
    .Y(_1715_));
 sky130_fd_sc_hd__xnor2_1 _4338_ (.A(_1699_),
    .B(_1715_),
    .Y(_1716_));
 sky130_fd_sc_hd__buf_2 _4339_ (.A(_1712_),
    .X(_1717_));
 sky130_fd_sc_hd__buf_2 _4340_ (.A(_1717_),
    .X(_1718_));
 sky130_fd_sc_hd__a22o_1 _4341_ (.A1(\sum[29] ),
    .A2(_1714_),
    .B1(_1716_),
    .B2(_1718_),
    .X(_0286_));
 sky130_fd_sc_hd__xor2_1 _4342_ (.A(_1697_),
    .B(_1698_),
    .X(_1719_));
 sky130_fd_sc_hd__a22o_1 _4343_ (.A1(\sum[28] ),
    .A2(_1714_),
    .B1(_1719_),
    .B2(_1718_),
    .X(_0285_));
 sky130_fd_sc_hd__a21oi_1 _4344_ (.A1(\sum[26] ),
    .A2(_1704_),
    .B1(_1695_),
    .Y(_1720_));
 sky130_fd_sc_hd__xnor2_1 _4345_ (.A(_1615_),
    .B(_1720_),
    .Y(_1721_));
 sky130_fd_sc_hd__a22o_1 _4346_ (.A1(\sum[27] ),
    .A2(_1714_),
    .B1(_1721_),
    .B2(_1718_),
    .X(_0284_));
 sky130_fd_sc_hd__clkbuf_2 _4347_ (.A(_1597_),
    .X(_1722_));
 sky130_fd_sc_hd__and3_1 _4348_ (.A(_1694_),
    .B(_1692_),
    .C(_1693_),
    .X(_1723_));
 sky130_fd_sc_hd__o21ai_1 _4349_ (.A1(_1695_),
    .A2(_1723_),
    .B1(_1717_),
    .Y(_1724_));
 sky130_fd_sc_hd__o21a_1 _4350_ (.A1(\sum[26] ),
    .A2(_1722_),
    .B1(_1724_),
    .X(_0283_));
 sky130_fd_sc_hd__buf_2 _4351_ (.A(_1605_),
    .X(_1725_));
 sky130_fd_sc_hd__a21bo_1 _4352_ (.A1(\sum[24] ),
    .A2(_1725_),
    .B1_N(_1690_),
    .X(_1726_));
 sky130_fd_sc_hd__nor2_1 _4353_ (.A(_1691_),
    .B(_1726_),
    .Y(_1727_));
 sky130_fd_sc_hd__a21o_1 _4354_ (.A1(_1691_),
    .A2(_1726_),
    .B1(_1707_),
    .X(_1728_));
 sky130_fd_sc_hd__o22a_1 _4355_ (.A1(\sum[25] ),
    .A2(_1598_),
    .B1(_1727_),
    .B2(_1728_),
    .X(_0282_));
 sky130_fd_sc_hd__buf_2 _4356_ (.A(_1717_),
    .X(_1729_));
 sky130_fd_sc_hd__or3_1 _4357_ (.A(_1685_),
    .B(_1688_),
    .C(_1689_),
    .X(_1730_));
 sky130_fd_sc_hd__a32o_1 _4358_ (.A1(_1729_),
    .A2(_1690_),
    .A3(_1730_),
    .B1(_1713_),
    .B2(\sum[24] ),
    .X(_0281_));
 sky130_fd_sc_hd__inv_2 _4359_ (.A(_1680_),
    .Y(_1731_));
 sky130_fd_sc_hd__nor2_1 _4360_ (.A(_1676_),
    .B(_1677_),
    .Y(_1732_));
 sky130_fd_sc_hd__o22a_1 _4361_ (.A1(\sum[21] ),
    .A2(_1614_),
    .B1(_1732_),
    .B2(_1686_),
    .X(_1733_));
 sky130_fd_sc_hd__and2_1 _4362_ (.A(_1731_),
    .B(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__o31a_1 _4363_ (.A1(_1678_),
    .A2(_1681_),
    .A3(_1734_),
    .B1(_1717_),
    .X(_1735_));
 sky130_fd_sc_hd__o21ai_1 _4364_ (.A1(_1678_),
    .A2(_1734_),
    .B1(_1681_),
    .Y(_1736_));
 sky130_fd_sc_hd__o2bb2a_1 _4365_ (.A1_N(_1735_),
    .A2_N(_1736_),
    .B1(_1722_),
    .B2(\sum[23] ),
    .X(_0280_));
 sky130_fd_sc_hd__nor2_1 _4366_ (.A(_1731_),
    .B(_1733_),
    .Y(_1737_));
 sky130_fd_sc_hd__nor2_1 _4367_ (.A(_1734_),
    .B(_1737_),
    .Y(_1738_));
 sky130_fd_sc_hd__o22a_1 _4368_ (.A1(\sum[22] ),
    .A2(_1722_),
    .B1(_1738_),
    .B2(_1711_),
    .X(_0279_));
 sky130_fd_sc_hd__buf_2 _4369_ (.A(_1597_),
    .X(_1739_));
 sky130_fd_sc_hd__a21o_1 _4370_ (.A1(\sum[20] ),
    .A2(_1704_),
    .B1(_1732_),
    .X(_1740_));
 sky130_fd_sc_hd__xnor2_1 _4371_ (.A(_1683_),
    .B(_1740_),
    .Y(_1741_));
 sky130_fd_sc_hd__o22a_1 _4372_ (.A1(\sum[21] ),
    .A2(_1739_),
    .B1(_1741_),
    .B2(_1711_),
    .X(_0278_));
 sky130_fd_sc_hd__buf_2 _4373_ (.A(_1713_),
    .X(_1742_));
 sky130_fd_sc_hd__nand2_1 _4374_ (.A(_1676_),
    .B(_1677_),
    .Y(_1743_));
 sky130_fd_sc_hd__nor2_1 _4375_ (.A(_1707_),
    .B(_1732_),
    .Y(_1744_));
 sky130_fd_sc_hd__a22o_1 _4376_ (.A1(\sum[20] ),
    .A2(_1742_),
    .B1(_1743_),
    .B2(_1744_),
    .X(_0277_));
 sky130_fd_sc_hd__nand2_1 _4377_ (.A(net378),
    .B(_1725_),
    .Y(_1745_));
 sky130_fd_sc_hd__nand2_1 _4378_ (.A(_1745_),
    .B(_1674_),
    .Y(_1746_));
 sky130_fd_sc_hd__o31a_1 _4379_ (.A1(_1669_),
    .A2(_1673_),
    .A3(_1746_),
    .B1(_1717_),
    .X(_1747_));
 sky130_fd_sc_hd__o21ai_1 _4380_ (.A1(_1669_),
    .A2(_1673_),
    .B1(_1746_),
    .Y(_1748_));
 sky130_fd_sc_hd__o2bb2a_1 _4381_ (.A1_N(_1747_),
    .A2_N(_1748_),
    .B1(_1722_),
    .B2(net378),
    .X(_0276_));
 sky130_fd_sc_hd__or2_1 _4382_ (.A(_1617_),
    .B(_1667_),
    .X(_1749_));
 sky130_fd_sc_hd__o21a_1 _4383_ (.A1(_1616_),
    .A2(_1749_),
    .B1(_1668_),
    .X(_1750_));
 sky130_fd_sc_hd__xnor2_1 _4384_ (.A(_1671_),
    .B(_1750_),
    .Y(_1751_));
 sky130_fd_sc_hd__o22a_1 _4385_ (.A1(\sum[18] ),
    .A2(_1598_),
    .B1(_1751_),
    .B2(_1711_),
    .X(_0275_));
 sky130_fd_sc_hd__nor2_1 _4386_ (.A(\sum[17] ),
    .B(_1704_),
    .Y(_1752_));
 sky130_fd_sc_hd__or2_1 _4387_ (.A(_1752_),
    .B(_1616_),
    .X(_1753_));
 sky130_fd_sc_hd__xnor2_1 _4388_ (.A(_1749_),
    .B(_1753_),
    .Y(_1754_));
 sky130_fd_sc_hd__o22a_1 _4389_ (.A1(\sum[17] ),
    .A2(_1739_),
    .B1(_1754_),
    .B2(_1708_),
    .X(_0274_));
 sky130_fd_sc_hd__dfrtp_1 _4390_ (.CLK(clknet_4_3_0_clock),
    .D(_0179_),
    .RESET_B(_0000_),
    .Q(\delta[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4391_ (.CLK(clknet_4_7_0_clock),
    .D(_0180_),
    .RESET_B(_0001_),
    .Q(net196));
 sky130_fd_sc_hd__dfrtp_1 _4392_ (.CLK(clknet_4_1_0_clock),
    .D(_0181_),
    .RESET_B(_0002_),
    .Q(net207));
 sky130_fd_sc_hd__dfrtp_1 _4393_ (.CLK(clknet_4_1_0_clock),
    .D(_0182_),
    .RESET_B(_0003_),
    .Q(net218));
 sky130_fd_sc_hd__dfrtp_1 _4394_ (.CLK(clknet_4_4_0_clock),
    .D(_0183_),
    .RESET_B(_0004_),
    .Q(net221));
 sky130_fd_sc_hd__dfrtp_1 _4395_ (.CLK(clknet_4_0_0_clock),
    .D(_0184_),
    .RESET_B(_0005_),
    .Q(net222));
 sky130_fd_sc_hd__dfrtp_1 _4396_ (.CLK(clknet_4_0_0_clock),
    .D(_0185_),
    .RESET_B(_0006_),
    .Q(net223));
 sky130_fd_sc_hd__dfrtp_1 _4397_ (.CLK(clknet_4_1_0_clock),
    .D(_0186_),
    .RESET_B(_0007_),
    .Q(net224));
 sky130_fd_sc_hd__dfrtp_1 _4398_ (.CLK(clknet_4_1_0_clock),
    .D(_0187_),
    .RESET_B(_0008_),
    .Q(net225));
 sky130_fd_sc_hd__dfrtp_1 _4399_ (.CLK(clknet_4_1_0_clock),
    .D(_0188_),
    .RESET_B(_0009_),
    .Q(net226));
 sky130_fd_sc_hd__dfrtp_1 _4400_ (.CLK(clknet_4_0_0_clock),
    .D(_0189_),
    .RESET_B(_0010_),
    .Q(net227));
 sky130_fd_sc_hd__dfrtp_1 _4401_ (.CLK(clknet_4_4_0_clock),
    .D(_0190_),
    .RESET_B(_0011_),
    .Q(net197));
 sky130_fd_sc_hd__dfrtp_1 _4402_ (.CLK(clknet_4_4_0_clock),
    .D(_0191_),
    .RESET_B(_0012_),
    .Q(net198));
 sky130_fd_sc_hd__dfrtp_1 _4403_ (.CLK(clknet_4_4_0_clock),
    .D(_0192_),
    .RESET_B(_0013_),
    .Q(net199));
 sky130_fd_sc_hd__dfrtp_1 _4404_ (.CLK(clknet_4_4_0_clock),
    .D(_0193_),
    .RESET_B(_0014_),
    .Q(net200));
 sky130_fd_sc_hd__dfrtp_1 _4405_ (.CLK(clknet_4_4_0_clock),
    .D(_0194_),
    .RESET_B(_0015_),
    .Q(net201));
 sky130_fd_sc_hd__dfrtp_1 _4406_ (.CLK(clknet_4_4_0_clock),
    .D(_0195_),
    .RESET_B(_0016_),
    .Q(net202));
 sky130_fd_sc_hd__dfrtp_1 _4407_ (.CLK(clknet_4_5_0_clock),
    .D(_0196_),
    .RESET_B(_0017_),
    .Q(net203));
 sky130_fd_sc_hd__dfrtp_1 _4408_ (.CLK(clknet_4_5_0_clock),
    .D(_0197_),
    .RESET_B(_0018_),
    .Q(net204));
 sky130_fd_sc_hd__dfrtp_1 _4409_ (.CLK(clknet_4_5_0_clock),
    .D(_0198_),
    .RESET_B(_0019_),
    .Q(net205));
 sky130_fd_sc_hd__dfrtp_1 _4410_ (.CLK(clknet_4_5_0_clock),
    .D(_0199_),
    .RESET_B(_0020_),
    .Q(net206));
 sky130_fd_sc_hd__dfrtp_1 _4411_ (.CLK(clknet_4_5_0_clock),
    .D(_0200_),
    .RESET_B(_0021_),
    .Q(net208));
 sky130_fd_sc_hd__dfrtp_1 _4412_ (.CLK(clknet_4_5_0_clock),
    .D(_0201_),
    .RESET_B(_0022_),
    .Q(net209));
 sky130_fd_sc_hd__dfrtp_1 _4413_ (.CLK(clknet_4_5_0_clock),
    .D(_0202_),
    .RESET_B(_0023_),
    .Q(net210));
 sky130_fd_sc_hd__dfrtp_1 _4414_ (.CLK(clknet_4_6_0_clock),
    .D(_0203_),
    .RESET_B(_0024_),
    .Q(net211));
 sky130_fd_sc_hd__dfrtp_1 _4415_ (.CLK(clknet_4_6_0_clock),
    .D(_0204_),
    .RESET_B(_0025_),
    .Q(net212));
 sky130_fd_sc_hd__dfrtp_1 _4416_ (.CLK(clknet_4_6_0_clock),
    .D(_0205_),
    .RESET_B(_0026_),
    .Q(net213));
 sky130_fd_sc_hd__dfrtp_1 _4417_ (.CLK(clknet_4_5_0_clock),
    .D(_0206_),
    .RESET_B(_0027_),
    .Q(net214));
 sky130_fd_sc_hd__dfrtp_1 _4418_ (.CLK(clknet_4_6_0_clock),
    .D(_0207_),
    .RESET_B(_0028_),
    .Q(net215));
 sky130_fd_sc_hd__dfrtp_1 _4419_ (.CLK(clknet_4_7_0_clock),
    .D(_0208_),
    .RESET_B(_0029_),
    .Q(net216));
 sky130_fd_sc_hd__dfrtp_1 _4420_ (.CLK(clknet_4_7_0_clock),
    .D(_0209_),
    .RESET_B(_0030_),
    .Q(net217));
 sky130_fd_sc_hd__dfrtp_1 _4421_ (.CLK(clknet_4_7_0_clock),
    .D(_0210_),
    .RESET_B(_0031_),
    .Q(net219));
 sky130_fd_sc_hd__dfrtp_1 _4422_ (.CLK(clknet_4_7_0_clock),
    .D(_0211_),
    .RESET_B(_0032_),
    .Q(net220));
 sky130_fd_sc_hd__dfrtp_2 _4423_ (.CLK(clknet_4_9_0_clock),
    .D(_0212_),
    .RESET_B(_0033_),
    .Q(net228));
 sky130_fd_sc_hd__dfrtp_1 _4424_ (.CLK(clknet_4_9_0_clock),
    .D(_0213_),
    .RESET_B(_0034_),
    .Q(net239));
 sky130_fd_sc_hd__dfrtp_1 _4425_ (.CLK(clknet_4_11_0_clock),
    .D(_0214_),
    .RESET_B(_0035_),
    .Q(net250));
 sky130_fd_sc_hd__dfrtp_1 _4426_ (.CLK(clknet_4_11_0_clock),
    .D(_0215_),
    .RESET_B(_0036_),
    .Q(net253));
 sky130_fd_sc_hd__dfrtp_2 _4427_ (.CLK(clknet_4_11_0_clock),
    .D(_0216_),
    .RESET_B(_0037_),
    .Q(net254));
 sky130_fd_sc_hd__dfrtp_1 _4428_ (.CLK(clknet_4_11_0_clock),
    .D(_0217_),
    .RESET_B(_0038_),
    .Q(net255));
 sky130_fd_sc_hd__dfrtp_1 _4429_ (.CLK(clknet_4_14_0_clock),
    .D(_0218_),
    .RESET_B(_0039_),
    .Q(net256));
 sky130_fd_sc_hd__dfrtp_1 _4430_ (.CLK(clknet_4_11_0_clock),
    .D(_0219_),
    .RESET_B(_0040_),
    .Q(net257));
 sky130_fd_sc_hd__dfrtp_1 _4431_ (.CLK(clknet_4_11_0_clock),
    .D(_0220_),
    .RESET_B(_0041_),
    .Q(net258));
 sky130_fd_sc_hd__dfrtp_1 _4432_ (.CLK(clknet_4_14_0_clock),
    .D(_0221_),
    .RESET_B(_0042_),
    .Q(net259));
 sky130_fd_sc_hd__dfrtp_1 _4433_ (.CLK(clknet_4_11_0_clock),
    .D(_0222_),
    .RESET_B(_0043_),
    .Q(net229));
 sky130_fd_sc_hd__dfrtp_1 _4434_ (.CLK(clknet_4_11_0_clock),
    .D(_0223_),
    .RESET_B(_0044_),
    .Q(net230));
 sky130_fd_sc_hd__dfrtp_1 _4435_ (.CLK(clknet_4_14_0_clock),
    .D(_0224_),
    .RESET_B(_0045_),
    .Q(net231));
 sky130_fd_sc_hd__dfrtp_1 _4436_ (.CLK(clknet_4_11_0_clock),
    .D(_0225_),
    .RESET_B(_0046_),
    .Q(net232));
 sky130_fd_sc_hd__dfrtp_1 _4437_ (.CLK(clknet_4_14_0_clock),
    .D(_0226_),
    .RESET_B(_0047_),
    .Q(net233));
 sky130_fd_sc_hd__dfrtp_1 _4438_ (.CLK(clknet_4_14_0_clock),
    .D(_0227_),
    .RESET_B(_0048_),
    .Q(net234));
 sky130_fd_sc_hd__dfrtp_1 _4439_ (.CLK(clknet_4_15_0_clock),
    .D(_0228_),
    .RESET_B(_0049_),
    .Q(net235));
 sky130_fd_sc_hd__dfrtp_1 _4440_ (.CLK(clknet_4_15_0_clock),
    .D(_0229_),
    .RESET_B(_0050_),
    .Q(net236));
 sky130_fd_sc_hd__dfrtp_1 _4441_ (.CLK(clknet_4_15_0_clock),
    .D(_0230_),
    .RESET_B(_0051_),
    .Q(net237));
 sky130_fd_sc_hd__dfrtp_1 _4442_ (.CLK(clknet_4_15_0_clock),
    .D(_0231_),
    .RESET_B(_0052_),
    .Q(net238));
 sky130_fd_sc_hd__dfrtp_1 _4443_ (.CLK(clknet_4_12_0_clock),
    .D(_0232_),
    .RESET_B(_0053_),
    .Q(net240));
 sky130_fd_sc_hd__dfrtp_1 _4444_ (.CLK(clknet_4_12_0_clock),
    .D(_0233_),
    .RESET_B(_0054_),
    .Q(net241));
 sky130_fd_sc_hd__dfrtp_1 _4445_ (.CLK(clknet_4_12_0_clock),
    .D(_0234_),
    .RESET_B(_0055_),
    .Q(net242));
 sky130_fd_sc_hd__dfrtp_1 _4446_ (.CLK(clknet_4_12_0_clock),
    .D(_0235_),
    .RESET_B(_0056_),
    .Q(net243));
 sky130_fd_sc_hd__dfrtp_1 _4447_ (.CLK(clknet_4_13_0_clock),
    .D(_0236_),
    .RESET_B(_0057_),
    .Q(net244));
 sky130_fd_sc_hd__dfrtp_1 _4448_ (.CLK(clknet_4_12_0_clock),
    .D(_0237_),
    .RESET_B(_0058_),
    .Q(net245));
 sky130_fd_sc_hd__dfrtp_1 _4449_ (.CLK(clknet_4_13_0_clock),
    .D(_0238_),
    .RESET_B(_0059_),
    .Q(net246));
 sky130_fd_sc_hd__dfrtp_1 _4450_ (.CLK(clknet_4_13_0_clock),
    .D(_0239_),
    .RESET_B(_0060_),
    .Q(net247));
 sky130_fd_sc_hd__dfrtp_1 _4451_ (.CLK(clknet_4_13_0_clock),
    .D(_0240_),
    .RESET_B(_0061_),
    .Q(net248));
 sky130_fd_sc_hd__dfrtp_1 _4452_ (.CLK(clknet_4_12_0_clock),
    .D(_0241_),
    .RESET_B(_0062_),
    .Q(net249));
 sky130_fd_sc_hd__dfrtp_1 _4453_ (.CLK(clknet_4_13_0_clock),
    .D(_0242_),
    .RESET_B(_0063_),
    .Q(net251));
 sky130_fd_sc_hd__dfrtp_1 _4454_ (.CLK(clknet_4_7_0_clock),
    .D(_0243_),
    .RESET_B(_0064_),
    .Q(net252));
 sky130_fd_sc_hd__dfrtp_1 _4455_ (.CLK(clknet_4_0_0_clock),
    .D(_0244_),
    .RESET_B(_0065_),
    .Q(net195));
 sky130_fd_sc_hd__dfrtp_1 _4456_ (.CLK(clknet_4_3_0_clock),
    .D(_0245_),
    .RESET_B(_0066_),
    .Q(while_flag));
 sky130_fd_sc_hd__dfrtp_1 _4457_ (.CLK(clknet_4_0_0_clock),
    .D(_0246_),
    .RESET_B(_0067_),
    .Q(modereg));
 sky130_fd_sc_hd__dfrtp_1 _4458_ (.CLK(clknet_4_2_0_clock),
    .D(_0247_),
    .RESET_B(_0068_),
    .Q(\selectslice[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4459_ (.CLK(clknet_4_2_0_clock),
    .D(_0248_),
    .RESET_B(_0069_),
    .Q(\selectslice[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4460_ (.CLK(clknet_4_3_0_clock),
    .D(_0249_),
    .RESET_B(_0070_),
    .Q(\x[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4461_ (.CLK(clknet_4_3_0_clock),
    .D(_0250_),
    .RESET_B(_0071_),
    .Q(\x[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4462_ (.CLK(clknet_4_3_0_clock),
    .D(_0251_),
    .RESET_B(_0072_),
    .Q(\x[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4463_ (.CLK(clknet_4_9_0_clock),
    .D(_0252_),
    .RESET_B(_0073_),
    .Q(\x[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4464_ (.CLK(clknet_4_3_0_clock),
    .D(_0253_),
    .RESET_B(_0074_),
    .Q(\x[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4465_ (.CLK(clknet_4_9_0_clock),
    .D(_0254_),
    .RESET_B(_0075_),
    .Q(\x[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4466_ (.CLK(clknet_4_9_0_clock),
    .D(_0255_),
    .RESET_B(_0076_),
    .Q(\x[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4467_ (.CLK(clknet_4_9_0_clock),
    .D(_0256_),
    .RESET_B(_0077_),
    .Q(\x[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4468_ (.CLK(clknet_4_2_0_clock),
    .D(_0257_),
    .RESET_B(_0078_),
    .Q(\sum[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4469_ (.CLK(clknet_4_2_0_clock),
    .D(_0258_),
    .RESET_B(_0079_),
    .Q(\sum[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4470_ (.CLK(clknet_4_0_0_clock),
    .D(_0259_),
    .RESET_B(_0080_),
    .Q(\sum[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4471_ (.CLK(clknet_4_2_0_clock),
    .D(_0260_),
    .RESET_B(_0081_),
    .Q(\sum[3] ));
 sky130_fd_sc_hd__dfrtp_4 _4472_ (.CLK(clknet_4_2_0_clock),
    .D(_0261_),
    .RESET_B(_0082_),
    .Q(\sum[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4473_ (.CLK(clknet_4_0_0_clock),
    .D(_0262_),
    .RESET_B(_0083_),
    .Q(\sum[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4474_ (.CLK(clknet_4_2_0_clock),
    .D(_0263_),
    .RESET_B(_0084_),
    .Q(\sum[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4475_ (.CLK(clknet_4_2_0_clock),
    .D(_0264_),
    .RESET_B(_0085_),
    .Q(\sum[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4476_ (.CLK(clknet_4_2_0_clock),
    .D(_0265_),
    .RESET_B(_0086_),
    .Q(\sum[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4477_ (.CLK(clknet_4_2_0_clock),
    .D(_0266_),
    .RESET_B(_0087_),
    .Q(\sum[9] ));
 sky130_fd_sc_hd__dfrtp_1 _4478_ (.CLK(clknet_4_2_0_clock),
    .D(_0267_),
    .RESET_B(_0088_),
    .Q(\sum[10] ));
 sky130_fd_sc_hd__dfrtp_1 _4479_ (.CLK(clknet_4_2_0_clock),
    .D(_0268_),
    .RESET_B(_0089_),
    .Q(\sum[11] ));
 sky130_fd_sc_hd__dfrtp_1 _4480_ (.CLK(clknet_4_2_0_clock),
    .D(_0269_),
    .RESET_B(_0090_),
    .Q(\sum[12] ));
 sky130_fd_sc_hd__dfrtp_1 _4481_ (.CLK(clknet_4_8_0_clock),
    .D(_0270_),
    .RESET_B(_0091_),
    .Q(\sum[13] ));
 sky130_fd_sc_hd__dfrtp_1 _4482_ (.CLK(clknet_4_2_0_clock),
    .D(_0271_),
    .RESET_B(_0092_),
    .Q(\sum[14] ));
 sky130_fd_sc_hd__dfrtp_1 _4483_ (.CLK(clknet_4_8_0_clock),
    .D(_0272_),
    .RESET_B(_0093_),
    .Q(\sum[15] ));
 sky130_fd_sc_hd__dfrtp_1 _4484_ (.CLK(clknet_4_9_0_clock),
    .D(_0273_),
    .RESET_B(_0094_),
    .Q(\sum[16] ));
 sky130_fd_sc_hd__dfrtp_1 _4485_ (.CLK(clknet_4_8_0_clock),
    .D(_0274_),
    .RESET_B(_0095_),
    .Q(\sum[17] ));
 sky130_fd_sc_hd__dfrtp_1 _4486_ (.CLK(clknet_4_9_0_clock),
    .D(_0275_),
    .RESET_B(_0096_),
    .Q(\sum[18] ));
 sky130_fd_sc_hd__dfrtp_1 _4487_ (.CLK(clknet_4_8_0_clock),
    .D(_0276_),
    .RESET_B(_0097_),
    .Q(\sum[19] ));
 sky130_fd_sc_hd__dfrtp_2 _4488_ (.CLK(clknet_4_8_0_clock),
    .D(_0277_),
    .RESET_B(_0098_),
    .Q(\sum[20] ));
 sky130_fd_sc_hd__dfrtp_2 _4489_ (.CLK(clknet_4_8_0_clock),
    .D(_0278_),
    .RESET_B(_0099_),
    .Q(\sum[21] ));
 sky130_fd_sc_hd__dfrtp_2 _4490_ (.CLK(clknet_4_8_0_clock),
    .D(_0279_),
    .RESET_B(_0100_),
    .Q(\sum[22] ));
 sky130_fd_sc_hd__dfrtp_2 _4491_ (.CLK(clknet_4_8_0_clock),
    .D(_0280_),
    .RESET_B(_0101_),
    .Q(\sum[23] ));
 sky130_fd_sc_hd__dfrtp_2 _4492_ (.CLK(clknet_4_8_0_clock),
    .D(_0281_),
    .RESET_B(_0102_),
    .Q(\sum[24] ));
 sky130_fd_sc_hd__dfrtp_2 _4493_ (.CLK(clknet_4_8_0_clock),
    .D(_0282_),
    .RESET_B(_0103_),
    .Q(\sum[25] ));
 sky130_fd_sc_hd__dfrtp_2 _4494_ (.CLK(clknet_4_10_0_clock),
    .D(_0283_),
    .RESET_B(_0104_),
    .Q(\sum[26] ));
 sky130_fd_sc_hd__dfrtp_2 _4495_ (.CLK(clknet_4_10_0_clock),
    .D(_0284_),
    .RESET_B(_0105_),
    .Q(\sum[27] ));
 sky130_fd_sc_hd__dfrtp_4 _4496_ (.CLK(clknet_4_10_0_clock),
    .D(_0285_),
    .RESET_B(_0106_),
    .Q(\sum[28] ));
 sky130_fd_sc_hd__dfrtp_1 _4497_ (.CLK(clknet_4_10_0_clock),
    .D(_0286_),
    .RESET_B(_0107_),
    .Q(\sum[29] ));
 sky130_fd_sc_hd__dfrtp_1 _4498_ (.CLK(clknet_4_10_0_clock),
    .D(_0287_),
    .RESET_B(_0108_),
    .Q(\sum[30] ));
 sky130_fd_sc_hd__dfrtp_4 _4499_ (.CLK(clknet_4_10_0_clock),
    .D(_0288_),
    .RESET_B(_0109_),
    .Q(\sum[31] ));
 sky130_fd_sc_hd__dfrtp_2 _4500_ (.CLK(clknet_4_0_0_clock),
    .D(net557),
    .RESET_B(_0110_),
    .Q(\workunit1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4501_ (.CLK(clknet_4_1_0_clock),
    .D(net518),
    .RESET_B(_0111_),
    .Q(\workunit1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4502_ (.CLK(clknet_4_1_0_clock),
    .D(_0291_),
    .RESET_B(_0112_),
    .Q(\workunit1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4503_ (.CLK(clknet_4_1_0_clock),
    .D(_0292_),
    .RESET_B(_0113_),
    .Q(\workunit1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4504_ (.CLK(clknet_4_1_0_clock),
    .D(_0293_),
    .RESET_B(_0114_),
    .Q(\workunit1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4505_ (.CLK(clknet_4_0_0_clock),
    .D(_0294_),
    .RESET_B(_0115_),
    .Q(\workunit1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4506_ (.CLK(clknet_4_4_0_clock),
    .D(_0295_),
    .RESET_B(_0116_),
    .Q(\workunit1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4507_ (.CLK(clknet_4_4_0_clock),
    .D(_0296_),
    .RESET_B(_0117_),
    .Q(\workunit1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4508_ (.CLK(clknet_4_4_0_clock),
    .D(_0297_),
    .RESET_B(_0118_),
    .Q(\workunit1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4509_ (.CLK(clknet_4_5_0_clock),
    .D(_0298_),
    .RESET_B(_0119_),
    .Q(\workunit1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _4510_ (.CLK(clknet_4_4_0_clock),
    .D(_0299_),
    .RESET_B(_0120_),
    .Q(\workunit1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _4511_ (.CLK(clknet_4_4_0_clock),
    .D(_0300_),
    .RESET_B(_0121_),
    .Q(\workunit1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _4512_ (.CLK(clknet_4_4_0_clock),
    .D(_0301_),
    .RESET_B(_0122_),
    .Q(\workunit1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _4513_ (.CLK(clknet_4_4_0_clock),
    .D(_0302_),
    .RESET_B(_0123_),
    .Q(\workunit1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _4514_ (.CLK(clknet_4_5_0_clock),
    .D(_0303_),
    .RESET_B(_0124_),
    .Q(\workunit1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _4515_ (.CLK(clknet_4_4_0_clock),
    .D(_0304_),
    .RESET_B(_0125_),
    .Q(\workunit1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _4516_ (.CLK(clknet_4_5_0_clock),
    .D(_0305_),
    .RESET_B(_0126_),
    .Q(\workunit1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _4517_ (.CLK(clknet_4_5_0_clock),
    .D(_0306_),
    .RESET_B(_0127_),
    .Q(\workunit1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _4518_ (.CLK(clknet_4_5_0_clock),
    .D(_0307_),
    .RESET_B(_0128_),
    .Q(\workunit1[18] ));
 sky130_fd_sc_hd__dfrtp_1 _4519_ (.CLK(clknet_4_6_0_clock),
    .D(_0308_),
    .RESET_B(_0129_),
    .Q(\workunit1[19] ));
 sky130_fd_sc_hd__dfrtp_1 _4520_ (.CLK(clknet_4_5_0_clock),
    .D(_0309_),
    .RESET_B(_0130_),
    .Q(\workunit1[20] ));
 sky130_fd_sc_hd__dfrtp_2 _4521_ (.CLK(clknet_4_4_0_clock),
    .D(_0310_),
    .RESET_B(_0131_),
    .Q(\workunit1[21] ));
 sky130_fd_sc_hd__dfrtp_1 _4522_ (.CLK(clknet_4_6_0_clock),
    .D(_0311_),
    .RESET_B(_0132_),
    .Q(\workunit1[22] ));
 sky130_fd_sc_hd__dfrtp_1 _4523_ (.CLK(clknet_4_6_0_clock),
    .D(_0312_),
    .RESET_B(_0133_),
    .Q(\workunit1[23] ));
 sky130_fd_sc_hd__dfrtp_1 _4524_ (.CLK(clknet_4_6_0_clock),
    .D(_0313_),
    .RESET_B(_0134_),
    .Q(\workunit1[24] ));
 sky130_fd_sc_hd__dfrtp_1 _4525_ (.CLK(clknet_4_7_0_clock),
    .D(_0314_),
    .RESET_B(_0135_),
    .Q(\workunit1[25] ));
 sky130_fd_sc_hd__dfrtp_1 _4526_ (.CLK(clknet_4_5_0_clock),
    .D(_0315_),
    .RESET_B(_0136_),
    .Q(\workunit1[26] ));
 sky130_fd_sc_hd__dfrtp_1 _4527_ (.CLK(clknet_4_6_0_clock),
    .D(_0316_),
    .RESET_B(_0137_),
    .Q(\workunit1[27] ));
 sky130_fd_sc_hd__dfrtp_1 _4528_ (.CLK(clknet_4_6_0_clock),
    .D(_0317_),
    .RESET_B(_0138_),
    .Q(\workunit1[28] ));
 sky130_fd_sc_hd__dfrtp_1 _4529_ (.CLK(clknet_4_6_0_clock),
    .D(_0318_),
    .RESET_B(_0139_),
    .Q(\workunit1[29] ));
 sky130_fd_sc_hd__dfrtp_1 _4530_ (.CLK(clknet_4_7_0_clock),
    .D(_0319_),
    .RESET_B(_0140_),
    .Q(\workunit1[30] ));
 sky130_fd_sc_hd__dfrtp_4 _4531_ (.CLK(clknet_4_7_0_clock),
    .D(_0320_),
    .RESET_B(_0141_),
    .Q(\workunit1[31] ));
 sky130_fd_sc_hd__dfrtp_1 _4532_ (.CLK(clknet_4_10_0_clock),
    .D(net578),
    .RESET_B(_0142_),
    .Q(\workunit2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4533_ (.CLK(clknet_4_10_0_clock),
    .D(net529),
    .RESET_B(_0143_),
    .Q(\workunit2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4534_ (.CLK(clknet_4_11_0_clock),
    .D(_0323_),
    .RESET_B(_0144_),
    .Q(\workunit2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4535_ (.CLK(clknet_4_11_0_clock),
    .D(_0324_),
    .RESET_B(_0145_),
    .Q(\workunit2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4536_ (.CLK(clknet_4_11_0_clock),
    .D(_0325_),
    .RESET_B(_0146_),
    .Q(\workunit2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4537_ (.CLK(clknet_4_14_0_clock),
    .D(_0326_),
    .RESET_B(_0147_),
    .Q(\workunit2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4538_ (.CLK(clknet_4_14_0_clock),
    .D(_0327_),
    .RESET_B(_0148_),
    .Q(\workunit2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4539_ (.CLK(clknet_4_14_0_clock),
    .D(_0328_),
    .RESET_B(_0149_),
    .Q(\workunit2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4540_ (.CLK(clknet_4_14_0_clock),
    .D(_0329_),
    .RESET_B(_0150_),
    .Q(\workunit2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4541_ (.CLK(clknet_4_14_0_clock),
    .D(_0330_),
    .RESET_B(_0151_),
    .Q(\workunit2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _4542_ (.CLK(clknet_4_14_0_clock),
    .D(_0331_),
    .RESET_B(_0152_),
    .Q(\workunit2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _4543_ (.CLK(clknet_4_15_0_clock),
    .D(_0332_),
    .RESET_B(_0153_),
    .Q(\workunit2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _4544_ (.CLK(clknet_4_14_0_clock),
    .D(_0333_),
    .RESET_B(_0154_),
    .Q(\workunit2[12] ));
 sky130_fd_sc_hd__dfrtp_1 _4545_ (.CLK(clknet_4_15_0_clock),
    .D(_0334_),
    .RESET_B(_0155_),
    .Q(\workunit2[13] ));
 sky130_fd_sc_hd__dfrtp_1 _4546_ (.CLK(clknet_4_15_0_clock),
    .D(_0335_),
    .RESET_B(_0156_),
    .Q(\workunit2[14] ));
 sky130_fd_sc_hd__dfrtp_1 _4547_ (.CLK(clknet_4_13_0_clock),
    .D(_0336_),
    .RESET_B(_0157_),
    .Q(\workunit2[15] ));
 sky130_fd_sc_hd__dfrtp_1 _4548_ (.CLK(clknet_4_13_0_clock),
    .D(_0337_),
    .RESET_B(_0158_),
    .Q(\workunit2[16] ));
 sky130_fd_sc_hd__dfrtp_1 _4549_ (.CLK(clknet_4_12_0_clock),
    .D(_0338_),
    .RESET_B(_0159_),
    .Q(\workunit2[17] ));
 sky130_fd_sc_hd__dfrtp_1 _4550_ (.CLK(clknet_4_12_0_clock),
    .D(_0339_),
    .RESET_B(_0160_),
    .Q(\workunit2[18] ));
 sky130_fd_sc_hd__dfrtp_1 _4551_ (.CLK(clknet_4_12_0_clock),
    .D(_0340_),
    .RESET_B(_0161_),
    .Q(\workunit2[19] ));
 sky130_fd_sc_hd__dfrtp_1 _4552_ (.CLK(clknet_4_12_0_clock),
    .D(_0341_),
    .RESET_B(_0162_),
    .Q(\workunit2[20] ));
 sky130_fd_sc_hd__dfrtp_1 _4553_ (.CLK(clknet_4_15_0_clock),
    .D(_0342_),
    .RESET_B(_0163_),
    .Q(\workunit2[21] ));
 sky130_fd_sc_hd__dfrtp_1 _4554_ (.CLK(clknet_4_12_0_clock),
    .D(_0343_),
    .RESET_B(_0164_),
    .Q(\workunit2[22] ));
 sky130_fd_sc_hd__dfrtp_1 _4555_ (.CLK(clknet_4_12_0_clock),
    .D(_0344_),
    .RESET_B(_0165_),
    .Q(\workunit2[23] ));
 sky130_fd_sc_hd__dfrtp_1 _4556_ (.CLK(clknet_4_13_0_clock),
    .D(_0345_),
    .RESET_B(_0166_),
    .Q(\workunit2[24] ));
 sky130_fd_sc_hd__dfrtp_1 _4557_ (.CLK(clknet_4_13_0_clock),
    .D(_0346_),
    .RESET_B(_0167_),
    .Q(\workunit2[25] ));
 sky130_fd_sc_hd__dfrtp_1 _4558_ (.CLK(clknet_4_13_0_clock),
    .D(_0347_),
    .RESET_B(_0168_),
    .Q(\workunit2[26] ));
 sky130_fd_sc_hd__dfrtp_1 _4559_ (.CLK(clknet_4_13_0_clock),
    .D(_0348_),
    .RESET_B(_0169_),
    .Q(\workunit2[27] ));
 sky130_fd_sc_hd__dfrtp_1 _4560_ (.CLK(clknet_4_13_0_clock),
    .D(_0349_),
    .RESET_B(_0170_),
    .Q(\workunit2[28] ));
 sky130_fd_sc_hd__dfrtp_1 _4561_ (.CLK(clknet_4_12_0_clock),
    .D(net511),
    .RESET_B(_0171_),
    .Q(\workunit2[29] ));
 sky130_fd_sc_hd__dfrtp_1 _4562_ (.CLK(clknet_4_13_0_clock),
    .D(_0351_),
    .RESET_B(_0172_),
    .Q(\workunit2[30] ));
 sky130_fd_sc_hd__dfrtp_4 _4563_ (.CLK(clknet_4_13_0_clock),
    .D(net484),
    .RESET_B(_0173_),
    .Q(\workunit2[31] ));
 sky130_fd_sc_hd__dfrtp_2 _4564_ (.CLK(clknet_4_3_0_clock),
    .D(_2190_),
    .RESET_B(_0174_),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4565_ (.CLK(clknet_4_3_0_clock),
    .D(_2191_),
    .RESET_B(_0175_),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4566_ (.CLK(clknet_4_3_0_clock),
    .D(_2192_),
    .RESET_B(_0176_),
    .Q(\state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4567_ (.CLK(clknet_4_3_0_clock),
    .D(_2193_),
    .RESET_B(_0177_),
    .Q(\state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4568_ (.CLK(clknet_4_3_0_clock),
    .D(_2194_),
    .RESET_B(_0178_),
    .Q(\state[4] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_887 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(net554),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(net548),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(net560),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(net542),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(net566),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(net476),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(net478),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(net460),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(net452),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(net474),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(net538),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(net516),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(net458),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(net558),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(net466),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(net544),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(net514),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(net497),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(net456),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(net568),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(net540),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(net562),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(net450),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(net487),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(net530),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(net454),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(net546),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(net552),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(net493),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(net448),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(net503),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(net536),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(net576),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(net574),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(net462),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(net581),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(net519),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(net468),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(net470),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(net507),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(net572),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(net512),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(net495),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(net527),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(net480),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(net564),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(net485),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(net499),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(net550),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(net491),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(net464),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(net472),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(net521),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(net509),
    .X(net54));
 sky130_fd_sc_hd__dlymetal6s2s_1 input55 (.A(net583),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(net489),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(net482),
    .X(net57));
 sky130_fd_sc_hd__dlymetal6s2s_1 input58 (.A(net579),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(net523),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(net505),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(net534),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(net525),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(net570),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(net501),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(key_in[0]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(key_in[100]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(key_in[101]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(key_in[102]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(key_in[103]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(key_in[104]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(key_in[105]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(key_in[106]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(key_in[107]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(key_in[108]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(key_in[109]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(key_in[10]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(key_in[110]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(key_in[111]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(key_in[112]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input80 (.A(key_in[113]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(key_in[114]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(key_in[115]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(key_in[116]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(key_in[117]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(key_in[118]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(key_in[119]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(key_in[11]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(key_in[120]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(key_in[121]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(key_in[122]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(key_in[123]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(key_in[124]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(key_in[125]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(key_in[126]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(key_in[127]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(key_in[12]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(key_in[13]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(key_in[14]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(key_in[15]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(key_in[16]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(key_in[17]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(key_in[18]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(key_in[19]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(key_in[1]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(key_in[20]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(key_in[21]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(key_in[22]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 input108 (.A(key_in[23]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(key_in[24]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 input110 (.A(key_in[25]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(key_in[26]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(key_in[27]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(key_in[28]),
    .X(net113));
 sky130_fd_sc_hd__buf_1 input114 (.A(key_in[29]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(key_in[2]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(key_in[30]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 input117 (.A(key_in[31]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(key_in[32]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(key_in[33]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(key_in[34]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 input121 (.A(key_in[35]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(key_in[36]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(key_in[37]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(key_in[38]),
    .X(net124));
 sky130_fd_sc_hd__buf_1 input125 (.A(key_in[39]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(key_in[3]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(key_in[40]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(key_in[41]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 input129 (.A(key_in[42]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(key_in[43]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(key_in[44]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(key_in[45]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(key_in[46]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(key_in[47]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(key_in[48]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(key_in[49]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(key_in[4]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(key_in[50]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(key_in[51]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(key_in[52]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 input141 (.A(key_in[53]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 input142 (.A(key_in[54]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(key_in[55]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(key_in[56]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 input145 (.A(key_in[57]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 input146 (.A(key_in[58]),
    .X(net146));
 sky130_fd_sc_hd__dlymetal6s2s_1 input147 (.A(key_in[59]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(key_in[5]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 input149 (.A(key_in[60]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 input150 (.A(key_in[61]),
    .X(net150));
 sky130_fd_sc_hd__buf_1 input151 (.A(key_in[62]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(key_in[63]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 input153 (.A(key_in[64]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 input154 (.A(key_in[65]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 input155 (.A(key_in[66]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 input156 (.A(key_in[67]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 input157 (.A(key_in[68]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 input158 (.A(key_in[69]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 input159 (.A(key_in[6]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 input160 (.A(key_in[70]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 input161 (.A(key_in[71]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 input162 (.A(key_in[72]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 input163 (.A(key_in[73]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(key_in[74]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 input165 (.A(key_in[75]),
    .X(net165));
 sky130_fd_sc_hd__buf_1 input166 (.A(key_in[76]),
    .X(net166));
 sky130_fd_sc_hd__buf_1 input167 (.A(key_in[77]),
    .X(net167));
 sky130_fd_sc_hd__buf_1 input168 (.A(key_in[78]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 input169 (.A(key_in[79]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 input170 (.A(key_in[7]),
    .X(net170));
 sky130_fd_sc_hd__buf_1 input171 (.A(key_in[80]),
    .X(net171));
 sky130_fd_sc_hd__buf_1 input172 (.A(key_in[81]),
    .X(net172));
 sky130_fd_sc_hd__buf_1 input173 (.A(key_in[82]),
    .X(net173));
 sky130_fd_sc_hd__buf_1 input174 (.A(key_in[83]),
    .X(net174));
 sky130_fd_sc_hd__buf_1 input175 (.A(key_in[84]),
    .X(net175));
 sky130_fd_sc_hd__buf_1 input176 (.A(key_in[85]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 input177 (.A(key_in[86]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 input178 (.A(key_in[87]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 input179 (.A(key_in[88]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 input180 (.A(key_in[89]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 input181 (.A(key_in[8]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_2 input182 (.A(key_in[90]),
    .X(net182));
 sky130_fd_sc_hd__dlymetal6s2s_1 input183 (.A(key_in[91]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_2 input184 (.A(key_in[92]),
    .X(net184));
 sky130_fd_sc_hd__dlymetal6s2s_1 input185 (.A(key_in[93]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 input186 (.A(key_in[94]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_2 input187 (.A(key_in[95]),
    .X(net187));
 sky130_fd_sc_hd__buf_1 input188 (.A(key_in[96]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 input189 (.A(key_in[97]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 input190 (.A(key_in[98]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 input191 (.A(key_in[99]),
    .X(net191));
 sky130_fd_sc_hd__buf_1 input192 (.A(key_in[9]),
    .X(net192));
 sky130_fd_sc_hd__buf_1 input193 (.A(net532),
    .X(net193));
 sky130_fd_sc_hd__dlymetal6s2s_1 input194 (.A(net446),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_4 output195 (.A(net195),
    .X(all_done));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(data_out1[0]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(data_out1[10]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(data_out1[11]));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(data_out1[12]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(data_out1[13]));
 sky130_fd_sc_hd__buf_2 output201 (.A(net201),
    .X(data_out1[14]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(data_out1[15]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net203),
    .X(data_out1[16]));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(data_out1[17]));
 sky130_fd_sc_hd__buf_2 output205 (.A(net205),
    .X(data_out1[18]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(data_out1[19]));
 sky130_fd_sc_hd__buf_2 output207 (.A(net207),
    .X(data_out1[1]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net208),
    .X(data_out1[20]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net209),
    .X(data_out1[21]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net210),
    .X(data_out1[22]));
 sky130_fd_sc_hd__buf_2 output211 (.A(net211),
    .X(data_out1[23]));
 sky130_fd_sc_hd__buf_2 output212 (.A(net212),
    .X(data_out1[24]));
 sky130_fd_sc_hd__buf_2 output213 (.A(net213),
    .X(data_out1[25]));
 sky130_fd_sc_hd__buf_2 output214 (.A(net214),
    .X(data_out1[26]));
 sky130_fd_sc_hd__buf_2 output215 (.A(net215),
    .X(data_out1[27]));
 sky130_fd_sc_hd__buf_2 output216 (.A(net216),
    .X(data_out1[28]));
 sky130_fd_sc_hd__buf_2 output217 (.A(net217),
    .X(data_out1[29]));
 sky130_fd_sc_hd__buf_2 output218 (.A(net218),
    .X(data_out1[2]));
 sky130_fd_sc_hd__buf_2 output219 (.A(net219),
    .X(data_out1[30]));
 sky130_fd_sc_hd__buf_2 output220 (.A(net220),
    .X(data_out1[31]));
 sky130_fd_sc_hd__buf_2 output221 (.A(net221),
    .X(data_out1[3]));
 sky130_fd_sc_hd__buf_2 output222 (.A(net222),
    .X(data_out1[4]));
 sky130_fd_sc_hd__buf_2 output223 (.A(net223),
    .X(data_out1[5]));
 sky130_fd_sc_hd__buf_2 output224 (.A(net224),
    .X(data_out1[6]));
 sky130_fd_sc_hd__buf_2 output225 (.A(net225),
    .X(data_out1[7]));
 sky130_fd_sc_hd__buf_2 output226 (.A(net226),
    .X(data_out1[8]));
 sky130_fd_sc_hd__buf_2 output227 (.A(net227),
    .X(data_out1[9]));
 sky130_fd_sc_hd__clkbuf_4 output228 (.A(net228),
    .X(data_out2[0]));
 sky130_fd_sc_hd__clkbuf_4 output229 (.A(net229),
    .X(data_out2[10]));
 sky130_fd_sc_hd__clkbuf_4 output230 (.A(net230),
    .X(data_out2[11]));
 sky130_fd_sc_hd__clkbuf_4 output231 (.A(net231),
    .X(data_out2[12]));
 sky130_fd_sc_hd__clkbuf_4 output232 (.A(net232),
    .X(data_out2[13]));
 sky130_fd_sc_hd__clkbuf_4 output233 (.A(net233),
    .X(data_out2[14]));
 sky130_fd_sc_hd__clkbuf_4 output234 (.A(net234),
    .X(data_out2[15]));
 sky130_fd_sc_hd__clkbuf_4 output235 (.A(net235),
    .X(data_out2[16]));
 sky130_fd_sc_hd__clkbuf_4 output236 (.A(net236),
    .X(data_out2[17]));
 sky130_fd_sc_hd__clkbuf_4 output237 (.A(net237),
    .X(data_out2[18]));
 sky130_fd_sc_hd__clkbuf_4 output238 (.A(net238),
    .X(data_out2[19]));
 sky130_fd_sc_hd__buf_2 output239 (.A(net239),
    .X(data_out2[1]));
 sky130_fd_sc_hd__clkbuf_4 output240 (.A(net240),
    .X(data_out2[20]));
 sky130_fd_sc_hd__clkbuf_4 output241 (.A(net241),
    .X(data_out2[21]));
 sky130_fd_sc_hd__clkbuf_4 output242 (.A(net242),
    .X(data_out2[22]));
 sky130_fd_sc_hd__buf_2 output243 (.A(net243),
    .X(data_out2[23]));
 sky130_fd_sc_hd__buf_2 output244 (.A(net244),
    .X(data_out2[24]));
 sky130_fd_sc_hd__buf_2 output245 (.A(net245),
    .X(data_out2[25]));
 sky130_fd_sc_hd__buf_2 output246 (.A(net246),
    .X(data_out2[26]));
 sky130_fd_sc_hd__buf_2 output247 (.A(net247),
    .X(data_out2[27]));
 sky130_fd_sc_hd__buf_2 output248 (.A(net248),
    .X(data_out2[28]));
 sky130_fd_sc_hd__buf_2 output249 (.A(net249),
    .X(data_out2[29]));
 sky130_fd_sc_hd__clkbuf_4 output250 (.A(net250),
    .X(data_out2[2]));
 sky130_fd_sc_hd__buf_2 output251 (.A(net251),
    .X(data_out2[30]));
 sky130_fd_sc_hd__buf_2 output252 (.A(net252),
    .X(data_out2[31]));
 sky130_fd_sc_hd__clkbuf_4 output253 (.A(net253),
    .X(data_out2[3]));
 sky130_fd_sc_hd__clkbuf_4 output254 (.A(net254),
    .X(data_out2[4]));
 sky130_fd_sc_hd__clkbuf_4 output255 (.A(net255),
    .X(data_out2[5]));
 sky130_fd_sc_hd__clkbuf_4 output256 (.A(net256),
    .X(data_out2[6]));
 sky130_fd_sc_hd__clkbuf_4 output257 (.A(net257),
    .X(data_out2[7]));
 sky130_fd_sc_hd__clkbuf_4 output258 (.A(net258),
    .X(data_out2[8]));
 sky130_fd_sc_hd__clkbuf_4 output259 (.A(net259),
    .X(data_out2[9]));
 sky130_fd_sc_hd__clkbuf_1 max_cap260 (.A(_0841_),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_2 fanout261 (.A(\state[3] ),
    .X(net261));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout262 (.A(\state[2] ),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_2 fanout263 (.A(\state[2] ),
    .X(net263));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout264 (.A(net265),
    .X(net264));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout265 (.A(\state[1] ),
    .X(net265));
 sky130_fd_sc_hd__buf_1 fanout266 (.A(\workunit2[30] ),
    .X(net266));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout267 (.A(\workunit2[29] ),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_2 fanout268 (.A(\workunit2[28] ),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_2 fanout269 (.A(\workunit2[27] ),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_2 fanout270 (.A(\workunit2[27] ),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_2 fanout271 (.A(\workunit2[26] ),
    .X(net271));
 sky130_fd_sc_hd__buf_1 fanout272 (.A(\workunit2[26] ),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_2 fanout273 (.A(net274),
    .X(net273));
 sky130_fd_sc_hd__buf_1 fanout274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout275 (.A(\workunit2[25] ),
    .X(net275));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout277 (.A(\workunit2[24] ),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_2 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_2 fanout279 (.A(\workunit2[23] ),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_2 fanout280 (.A(\workunit2[22] ),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_2 fanout281 (.A(\workunit2[22] ),
    .X(net281));
 sky130_fd_sc_hd__buf_2 fanout282 (.A(\workunit2[21] ),
    .X(net282));
 sky130_fd_sc_hd__buf_1 fanout283 (.A(\workunit2[21] ),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_2 fanout284 (.A(\workunit2[20] ),
    .X(net284));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout285 (.A(\workunit2[20] ),
    .X(net285));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout286 (.A(net288),
    .X(net286));
 sky130_fd_sc_hd__buf_1 fanout287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout288 (.A(\workunit2[19] ),
    .X(net288));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout289 (.A(net290),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_2 fanout290 (.A(\workunit2[18] ),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_2 fanout291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout292 (.A(\workunit2[17] ),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_2 fanout293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout294 (.A(\workunit2[16] ),
    .X(net294));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__buf_1 fanout296 (.A(\workunit2[15] ),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_2 fanout297 (.A(net298),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_2 fanout298 (.A(\workunit2[14] ),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_2 fanout299 (.A(net300),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_2 fanout300 (.A(\workunit2[13] ),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_2 fanout301 (.A(net302),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_2 fanout302 (.A(\workunit2[12] ),
    .X(net302));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout303 (.A(net304),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_2 fanout304 (.A(\workunit2[11] ),
    .X(net304));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_2 fanout306 (.A(\workunit2[10] ),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_2 fanout307 (.A(net308),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_2 fanout308 (.A(\workunit2[9] ),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_2 fanout309 (.A(net310),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_2 fanout310 (.A(\workunit2[8] ),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_2 fanout311 (.A(\workunit2[7] ),
    .X(net311));
 sky130_fd_sc_hd__buf_1 fanout312 (.A(\workunit2[7] ),
    .X(net312));
 sky130_fd_sc_hd__buf_2 fanout313 (.A(\workunit2[6] ),
    .X(net313));
 sky130_fd_sc_hd__buf_1 fanout314 (.A(\workunit2[6] ),
    .X(net314));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout315 (.A(net316),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_2 fanout316 (.A(\workunit2[5] ),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_2 fanout317 (.A(\workunit2[4] ),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_2 fanout318 (.A(\workunit2[3] ),
    .X(net318));
 sky130_fd_sc_hd__buf_1 fanout319 (.A(net320),
    .X(net319));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout320 (.A(\workunit2[2] ),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_2 fanout321 (.A(\workunit2[1] ),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_2 fanout322 (.A(\workunit2[0] ),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_2 fanout323 (.A(\workunit1[30] ),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_2 fanout324 (.A(\workunit1[29] ),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_2 fanout325 (.A(\workunit1[28] ),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_2 fanout326 (.A(\workunit1[27] ),
    .X(net326));
 sky130_fd_sc_hd__buf_1 fanout327 (.A(\workunit1[27] ),
    .X(net327));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout328 (.A(net329),
    .X(net328));
 sky130_fd_sc_hd__buf_2 fanout329 (.A(\workunit1[26] ),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_2 fanout330 (.A(net331),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_2 fanout331 (.A(\workunit1[25] ),
    .X(net331));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout332 (.A(net333),
    .X(net332));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout333 (.A(\workunit1[24] ),
    .X(net333));
 sky130_fd_sc_hd__buf_2 fanout334 (.A(\workunit1[23] ),
    .X(net334));
 sky130_fd_sc_hd__buf_1 fanout335 (.A(\workunit1[23] ),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_2 fanout336 (.A(net337),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_2 fanout337 (.A(\workunit1[22] ),
    .X(net337));
 sky130_fd_sc_hd__buf_2 fanout338 (.A(\workunit1[21] ),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_2 fanout339 (.A(net340),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_2 fanout340 (.A(\workunit1[20] ),
    .X(net340));
 sky130_fd_sc_hd__buf_2 fanout341 (.A(net343),
    .X(net341));
 sky130_fd_sc_hd__buf_1 fanout342 (.A(net343),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 fanout343 (.A(\workunit1[19] ),
    .X(net343));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout344 (.A(net345),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_2 fanout345 (.A(\workunit1[18] ),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_2 fanout346 (.A(net347),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_2 fanout347 (.A(\workunit1[17] ),
    .X(net347));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout348 (.A(net349),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_2 fanout349 (.A(\workunit1[16] ),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_2 fanout350 (.A(net351),
    .X(net350));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout351 (.A(\workunit1[15] ),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_2 fanout352 (.A(net353),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_2 fanout353 (.A(\workunit1[14] ),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_2 fanout354 (.A(net355),
    .X(net354));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout355 (.A(\workunit1[13] ),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_2 fanout356 (.A(net357),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_2 fanout357 (.A(\workunit1[12] ),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_2 fanout358 (.A(\workunit1[11] ),
    .X(net358));
 sky130_fd_sc_hd__buf_1 fanout359 (.A(\workunit1[11] ),
    .X(net359));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout360 (.A(net361),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_2 fanout361 (.A(\workunit1[10] ),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_2 fanout362 (.A(net363),
    .X(net362));
 sky130_fd_sc_hd__buf_2 fanout363 (.A(\workunit1[9] ),
    .X(net363));
 sky130_fd_sc_hd__buf_2 fanout364 (.A(\workunit1[8] ),
    .X(net364));
 sky130_fd_sc_hd__buf_1 fanout365 (.A(\workunit1[8] ),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_2 fanout366 (.A(\workunit1[7] ),
    .X(net366));
 sky130_fd_sc_hd__buf_1 fanout367 (.A(\workunit1[7] ),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_2 fanout368 (.A(\workunit1[6] ),
    .X(net368));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout369 (.A(\workunit1[6] ),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_2 fanout370 (.A(net371),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_2 fanout371 (.A(\workunit1[5] ),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_2 fanout372 (.A(\workunit1[4] ),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_2 fanout373 (.A(\workunit1[3] ),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_2 fanout374 (.A(\workunit1[2] ),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_2 fanout375 (.A(\workunit1[1] ),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_2 fanout376 (.A(net377),
    .X(net376));
 sky130_fd_sc_hd__buf_1 fanout377 (.A(\workunit1[0] ),
    .X(net377));
 sky130_fd_sc_hd__buf_2 fanout378 (.A(\sum[19] ),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_2 fanout379 (.A(\sum[12] ),
    .X(net379));
 sky130_fd_sc_hd__buf_2 fanout380 (.A(net381),
    .X(net380));
 sky130_fd_sc_hd__buf_1 fanout381 (.A(\sum[11] ),
    .X(net381));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout382 (.A(\sum[9] ),
    .X(net382));
 sky130_fd_sc_hd__buf_2 fanout383 (.A(\sum[6] ),
    .X(net383));
 sky130_fd_sc_hd__buf_1 fanout384 (.A(\sum[1] ),
    .X(net384));
 sky130_fd_sc_hd__buf_2 fanout385 (.A(\sum[0] ),
    .X(net385));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout386 (.A(net387),
    .X(net386));
 sky130_fd_sc_hd__buf_1 fanout387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout388 (.A(net389),
    .X(net388));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout389 (.A(net391),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_2 fanout390 (.A(net391),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_2 fanout391 (.A(\selectslice[1] ),
    .X(net391));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout392 (.A(net393),
    .X(net392));
 sky130_fd_sc_hd__buf_1 fanout393 (.A(net394),
    .X(net393));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout394 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__buf_1 fanout395 (.A(net397),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_2 fanout396 (.A(net397),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_2 fanout397 (.A(\selectslice[0] ),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_2 fanout398 (.A(net399),
    .X(net398));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout399 (.A(\delta[0] ),
    .X(net399));
 sky130_fd_sc_hd__buf_2 fanout400 (.A(net401),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_2 fanout401 (.A(net404),
    .X(net401));
 sky130_fd_sc_hd__buf_2 fanout402 (.A(net403),
    .X(net402));
 sky130_fd_sc_hd__buf_2 fanout403 (.A(net404),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_2 fanout404 (.A(net421),
    .X(net404));
 sky130_fd_sc_hd__buf_2 fanout405 (.A(net409),
    .X(net405));
 sky130_fd_sc_hd__buf_2 fanout406 (.A(net409),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_4 fanout407 (.A(net409),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_2 fanout408 (.A(net409),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_2 fanout409 (.A(net421),
    .X(net409));
 sky130_fd_sc_hd__buf_2 fanout410 (.A(net413),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_4 fanout411 (.A(net413),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_2 fanout412 (.A(net413),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_2 fanout413 (.A(net420),
    .X(net413));
 sky130_fd_sc_hd__buf_2 fanout414 (.A(net418),
    .X(net414));
 sky130_fd_sc_hd__buf_2 fanout415 (.A(net417),
    .X(net415));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout416 (.A(net417),
    .X(net416));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__buf_1 fanout418 (.A(net420),
    .X(net418));
 sky130_fd_sc_hd__buf_2 fanout419 (.A(net420),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_2 fanout420 (.A(net421),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_2 fanout421 (.A(net447),
    .X(net421));
 sky130_fd_sc_hd__buf_2 fanout422 (.A(net423),
    .X(net422));
 sky130_fd_sc_hd__buf_1 fanout423 (.A(net434),
    .X(net423));
 sky130_fd_sc_hd__buf_2 fanout424 (.A(net426),
    .X(net424));
 sky130_fd_sc_hd__buf_2 fanout425 (.A(net426),
    .X(net425));
 sky130_fd_sc_hd__buf_1 fanout426 (.A(net434),
    .X(net426));
 sky130_fd_sc_hd__buf_2 fanout427 (.A(net429),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_2 fanout428 (.A(net429),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_2 fanout429 (.A(net432),
    .X(net429));
 sky130_fd_sc_hd__buf_2 fanout430 (.A(net432),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_2 fanout431 (.A(net432),
    .X(net431));
 sky130_fd_sc_hd__buf_1 fanout432 (.A(net433),
    .X(net432));
 sky130_fd_sc_hd__buf_2 fanout433 (.A(net434),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_2 fanout434 (.A(net445),
    .X(net434));
 sky130_fd_sc_hd__buf_2 fanout435 (.A(net436),
    .X(net435));
 sky130_fd_sc_hd__buf_2 fanout436 (.A(net439),
    .X(net436));
 sky130_fd_sc_hd__buf_2 fanout437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_2 fanout438 (.A(net439),
    .X(net438));
 sky130_fd_sc_hd__buf_1 fanout439 (.A(net445),
    .X(net439));
 sky130_fd_sc_hd__buf_2 fanout440 (.A(net443),
    .X(net440));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout441 (.A(net444),
    .X(net441));
 sky130_fd_sc_hd__buf_2 fanout442 (.A(net443),
    .X(net442));
 sky130_fd_sc_hd__buf_2 fanout443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__buf_2 fanout444 (.A(net445),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_2 fanout445 (.A(net447),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clock (.A(clock),
    .X(clknet_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clock (.A(clknet_0_clock),
    .X(clknet_4_0_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clock (.A(clknet_0_clock),
    .X(clknet_4_1_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clock (.A(clknet_0_clock),
    .X(clknet_4_2_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clock (.A(clknet_0_clock),
    .X(clknet_4_3_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clock (.A(clknet_0_clock),
    .X(clknet_4_4_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clock (.A(clknet_0_clock),
    .X(clknet_4_5_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clock (.A(clknet_0_clock),
    .X(clknet_4_6_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clock (.A(clknet_0_clock),
    .X(clknet_4_7_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clock (.A(clknet_0_clock),
    .X(clknet_4_8_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clock (.A(clknet_0_clock),
    .X(clknet_4_9_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clock (.A(clknet_0_clock),
    .X(clknet_4_10_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clock (.A(clknet_0_clock),
    .X(clknet_4_11_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clock (.A(clknet_0_clock),
    .X(clknet_4_12_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clock (.A(clknet_0_clock),
    .X(clknet_4_13_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clock (.A(clknet_0_clock),
    .X(clknet_4_14_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clock (.A(clknet_0_clock),
    .X(clknet_4_15_0_clock));
 sky130_fd_sc_hd__inv_6 clkload0 (.A(clknet_4_0_0_clock));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_4_1_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkload2 (.A(clknet_4_2_0_clock));
 sky130_fd_sc_hd__clkinvlp_4 clkload3 (.A(clknet_4_3_0_clock));
 sky130_fd_sc_hd__clkbuf_4 clkload4 (.A(clknet_4_5_0_clock));
 sky130_fd_sc_hd__clkinvlp_4 clkload5 (.A(clknet_4_6_0_clock));
 sky130_fd_sc_hd__inv_6 clkload6 (.A(clknet_4_7_0_clock));
 sky130_fd_sc_hd__clkinv_4 clkload7 (.A(clknet_4_8_0_clock));
 sky130_fd_sc_hd__inv_6 clkload8 (.A(clknet_4_9_0_clock));
 sky130_fd_sc_hd__inv_6 clkload9 (.A(clknet_4_10_0_clock));
 sky130_fd_sc_hd__bufinv_16 clkload10 (.A(clknet_4_11_0_clock));
 sky130_fd_sc_hd__clkinv_2 clkload11 (.A(clknet_4_12_0_clock));
 sky130_fd_sc_hd__clkbuf_8 clkload12 (.A(clknet_4_13_0_clock));
 sky130_fd_sc_hd__bufinv_16 clkload13 (.A(clknet_4_14_0_clock));
 sky130_fd_sc_hd__inv_6 clkload14 (.A(clknet_4_15_0_clock));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(reset),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net194),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(data_in1[7]),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net30),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(data_in1[2]),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net23),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(data_in1[17]),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net9),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(data_in1[3]),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net26),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(data_in1[26]),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net19),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(data_in1[20]),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net13),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(data_in1[16]),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net8),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(data_in2[11]),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net35),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(data_in2[26]),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net51),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(data_in1[22]),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net15),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(data_in2[14]),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net38),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(data_in2[15]),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net39),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(data_in2[27]),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net52),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(data_in1[18]),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net10),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(data_in1[14]),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net6),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(data_in1[15]),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net7),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(data_in2[20]),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net45),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(data_in2[31]),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net57),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_0352_),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(data_in2[22]),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net47),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(data_in1[30]),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net24),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(data_in2[30]),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net56),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(data_in2[25]),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net50),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(data_in1[6]),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net29),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(data_in2[19]),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net43),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(data_in1[25]),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net18),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(data_in2[23]),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net48),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(data_in2[9]),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net64),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(data_in1[8]),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net31),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(data_in2[5]),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net60),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(data_in2[16]),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net40),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(data_in2[29]),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net54),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0350_),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(data_in2[18]),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net42),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(data_in1[24]),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net17),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(data_in1[1]),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net12),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_0290_),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(data_in2[13]),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net37),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(data_in2[28]),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net53),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(data_in2[4]),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net59),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(data_in2[7]),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net62),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(data_in2[1]),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net44),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0322_),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(data_in1[31]),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net25),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(mode),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net193),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(data_in2[6]),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net61),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(data_in1[9]),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net32),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(data_in1[19]),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net11),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(data_in1[28]),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net21),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(data_in1[12]),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net4),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(data_in1[23]),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net16),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(data_in1[4]),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(net27),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(data_in1[10]),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net2),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(data_in2[24]),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(net49),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(data_in1[5]),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(net28),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(data_in1[0]),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(net1),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_1591_),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0289_),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(data_in1[21]),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(net14),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(data_in1[11]),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net3),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(data_in1[29]),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(net22),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(data_in2[21]),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(net46),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(data_in1[13]),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(net5),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(data_in1[27]),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(net20),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(data_in2[8]),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(net63),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(data_in2[17]),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(net41),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(data_in2[10]),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(net34),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(data_in2[0]),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(net33),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_0321_),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(data_in2[3]),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(net58),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(data_in2[12]),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(net36),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(data_in2[2]),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(net55),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\x[7] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\x[1] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\x[3] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\x[2] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\x[4] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\x[5] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\sum[1] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\sum[13] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\sum[3] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\sum[8] ),
    .X(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(data_in1[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(data_in2[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\workunit1[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_0874_));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_477 ();
endmodule
