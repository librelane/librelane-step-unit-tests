../002-success-flatten/spm.spice