../001-success/aes_example.lef