../001-success/spm.lef