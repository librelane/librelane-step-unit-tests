../001-success_explicit/dummy_doubleheight.lef