../../klayout.streamout/002-success_macros/user_proj_example2.lef