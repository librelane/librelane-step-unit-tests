VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spm
  CLASS BLOCK ;
  FOREIGN spm ;
  ORIGIN 0.000 0.000 ;
  SIZE 101.205 BY 111.925 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.280 20.380 95.920 21.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 15.020 10.640 16.620 100.880 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.280 17.080 95.920 18.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 11.720 10.640 13.320 100.880 ;
    END
  END VPWR
  PIN clk
    ANTENNAGATEAREA 10.176000 ;
    PORT
      LAYER met3 ;
        RECT 97.205 54.440 101.205 55.040 ;
    END
  END clk
  PIN p
    ANTENNAGATEAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END p
  PIN rst
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END rst
  PIN x[0]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 7.450 107.925 7.730 111.925 ;
    END
  END x[0]
  PIN x[10]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.050 107.925 35.330 111.925 ;
    END
  END x[10]
  PIN x[11]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 37.810 107.925 38.090 111.925 ;
    END
  END x[11]
  PIN x[12]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 40.570 107.925 40.850 111.925 ;
    END
  END x[12]
  PIN x[13]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 43.330 107.925 43.610 111.925 ;
    END
  END x[13]
  PIN x[14]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 46.090 107.925 46.370 111.925 ;
    END
  END x[14]
  PIN x[15]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 48.850 107.925 49.130 111.925 ;
    END
  END x[15]
  PIN x[16]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 107.925 51.890 111.925 ;
    END
  END x[16]
  PIN x[17]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.370 107.925 54.650 111.925 ;
    END
  END x[17]
  PIN x[18]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 57.130 107.925 57.410 111.925 ;
    END
  END x[18]
  PIN x[19]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 59.890 107.925 60.170 111.925 ;
    END
  END x[19]
  PIN x[1]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 10.210 107.925 10.490 111.925 ;
    END
  END x[1]
  PIN x[20]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 62.650 107.925 62.930 111.925 ;
    END
  END x[20]
  PIN x[21]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 65.410 107.925 65.690 111.925 ;
    END
  END x[21]
  PIN x[22]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 68.170 107.925 68.450 111.925 ;
    END
  END x[22]
  PIN x[23]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 107.925 71.210 111.925 ;
    END
  END x[23]
  PIN x[24]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 73.690 107.925 73.970 111.925 ;
    END
  END x[24]
  PIN x[25]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 76.450 107.925 76.730 111.925 ;
    END
  END x[25]
  PIN x[26]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 79.210 107.925 79.490 111.925 ;
    END
  END x[26]
  PIN x[27]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 81.970 107.925 82.250 111.925 ;
    END
  END x[27]
  PIN x[28]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 84.730 107.925 85.010 111.925 ;
    END
  END x[28]
  PIN x[29]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 87.490 107.925 87.770 111.925 ;
    END
  END x[29]
  PIN x[2]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 12.970 107.925 13.250 111.925 ;
    END
  END x[2]
  PIN x[30]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 107.925 90.530 111.925 ;
    END
  END x[30]
  PIN x[31]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 93.010 107.925 93.290 111.925 ;
    END
  END x[31]
  PIN x[3]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 15.730 107.925 16.010 111.925 ;
    END
  END x[3]
  PIN x[4]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 18.490 107.925 18.770 111.925 ;
    END
  END x[4]
  PIN x[5]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 21.250 107.925 21.530 111.925 ;
    END
  END x[5]
  PIN x[6]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 24.010 107.925 24.290 111.925 ;
    END
  END x[6]
  PIN x[7]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 26.770 107.925 27.050 111.925 ;
    END
  END x[7]
  PIN x[8]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.530 107.925 29.810 111.925 ;
    END
  END x[8]
  PIN x[9]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 107.925 32.570 111.925 ;
    END
  END x[9]
  PIN y
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END y
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 95.680 100.725 ;
      LAYER met1 ;
        RECT 4.670 10.640 95.680 100.880 ;
      LAYER met2 ;
        RECT 4.690 107.645 7.170 108.530 ;
        RECT 8.010 107.645 9.930 108.530 ;
        RECT 10.770 107.645 12.690 108.530 ;
        RECT 13.530 107.645 15.450 108.530 ;
        RECT 16.290 107.645 18.210 108.530 ;
        RECT 19.050 107.645 20.970 108.530 ;
        RECT 21.810 107.645 23.730 108.530 ;
        RECT 24.570 107.645 26.490 108.530 ;
        RECT 27.330 107.645 29.250 108.530 ;
        RECT 30.090 107.645 32.010 108.530 ;
        RECT 32.850 107.645 34.770 108.530 ;
        RECT 35.610 107.645 37.530 108.530 ;
        RECT 38.370 107.645 40.290 108.530 ;
        RECT 41.130 107.645 43.050 108.530 ;
        RECT 43.890 107.645 45.810 108.530 ;
        RECT 46.650 107.645 48.570 108.530 ;
        RECT 49.410 107.645 51.330 108.530 ;
        RECT 52.170 107.645 54.090 108.530 ;
        RECT 54.930 107.645 56.850 108.530 ;
        RECT 57.690 107.645 59.610 108.530 ;
        RECT 60.450 107.645 62.370 108.530 ;
        RECT 63.210 107.645 65.130 108.530 ;
        RECT 65.970 107.645 67.890 108.530 ;
        RECT 68.730 107.645 70.650 108.530 ;
        RECT 71.490 107.645 73.410 108.530 ;
        RECT 74.250 107.645 76.170 108.530 ;
        RECT 77.010 107.645 78.930 108.530 ;
        RECT 79.770 107.645 81.690 108.530 ;
        RECT 82.530 107.645 84.450 108.530 ;
        RECT 85.290 107.645 87.210 108.530 ;
        RECT 88.050 107.645 89.970 108.530 ;
        RECT 90.810 107.645 92.730 108.530 ;
        RECT 93.570 107.645 94.200 108.530 ;
        RECT 4.690 4.280 94.200 107.645 ;
        RECT 4.690 4.000 75.250 4.280 ;
        RECT 76.090 4.000 94.200 4.280 ;
      LAYER met3 ;
        RECT 4.000 84.000 97.205 100.805 ;
        RECT 4.400 82.600 97.205 84.000 ;
        RECT 4.000 55.440 97.205 82.600 ;
        RECT 4.000 54.040 96.805 55.440 ;
        RECT 4.000 28.240 97.205 54.040 ;
        RECT 4.400 26.840 97.205 28.240 ;
        RECT 4.000 10.715 97.205 26.840 ;
      LAYER met4 ;
        RECT 86.775 36.895 87.105 97.065 ;
  END
END spm
END LIBRARY

