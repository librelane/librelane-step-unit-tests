../../klayout.streamout/002-success_macros/user_proj_example.lef