module manual_macro_placement_test (clk1,
    clk2,
    p1,
    p2,
    rst1,
    rst2,
    y1,
    y2,
    x1,
    x2);
 input clk1;
 input clk2;
 output p1;
 output p2;
 input rst1;
 input rst2;
 input y1;
 input y2;
 input [31:0] x1;
 input [31:0] x2;

 wire tmp;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;

 sky130_fd_sc_hd__clkbuf_1 buffer (.A(tmp),
    .X(net70));
 spm spm_inst_0 (.clk(clk1),
    .p(net69),
    .rst(net1),
    .y(net67),
    .x({net27,
    net26,
    net24,
    net23,
    net22,
    net21,
    net20,
    net19,
    net18,
    net17,
    net16,
    net15,
    net13,
    net12,
    net11,
    net10,
    net9,
    net8,
    net7,
    net6,
    net5,
    net4,
    net34,
    net33,
    net32,
    net31,
    net30,
    net29,
    net28,
    net25,
    net14,
    net3}));
 spm spm_inst_1 (.clk(clk2),
    .p(tmp),
    .rst(net2),
    .y(net68),
    .x({net59,
    net58,
    net56,
    net55,
    net54,
    net53,
    net52,
    net51,
    net50,
    net49,
    net48,
    net47,
    net45,
    net44,
    net43,
    net42,
    net41,
    net40,
    net39,
    net38,
    net37,
    net36,
    net66,
    net65,
    net64,
    net63,
    net62,
    net61,
    net60,
    net57,
    net46,
    net35}));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Left_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Left_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Left_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Left_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Left_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Left_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Left_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Left_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Left_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Left_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Left_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Left_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Left_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Left_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Left_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Left_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Left_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Left_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Left_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Left_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Left_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Left_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Left_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Left_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Left_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Left_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Left_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_3_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_3_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_3_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_3_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_3_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_3_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_3_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_3_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_3_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_3_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_3_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_3_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_3_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_3_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_3_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_3_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_3_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_3_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_3_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_3_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_3_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_3_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_3_Right_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_3_Right_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_3_Right_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_3_Right_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_3_Right_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_3_Right_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_3_Right_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_3_Right_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_3_Right_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_3_Right_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_3_Right_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_3_Right_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_3_Right_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_3_Right_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_3_Right_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_3_Right_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_3_Right_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_3_Right_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_3_Right_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_3_Right_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_3_Right_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_3_Right_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_3_Right_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_3_Right_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_3_Right_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_3_Right_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_3_Right_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_3_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_3_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_3_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_3_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_3_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_3_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_3_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_3_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_3_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_3_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_3_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_3_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_3_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_3_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_3_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_3_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_3_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_3_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_3_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_3_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_3_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_3_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_3_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_3_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_3_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_3_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_3_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_3_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_3_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_3_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_3_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_3_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_3_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_3_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_3_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_3_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_3_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_3_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_3_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_3_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_3_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_3_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_3_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_3_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_3_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_3_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_3_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_3_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_3_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Right_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Right_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Right_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Right_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Right_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Right_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Right_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Right_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Right_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Right_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Right_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Right_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Right_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Right_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Right_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Right_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Right_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Right_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Right_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Right_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Right_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Right_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Right_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Right_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Right_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Right_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Right_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Right_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Right_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Right_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Right_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Right_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Right_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Right_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Right_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Right_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Right_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Right_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Right_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Right_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Right_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Right_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Right_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Right_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Right_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Right_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Right_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Right_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Right_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_3_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_3_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_3_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_3_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_3_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_3_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_3_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_3_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_3_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_3_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_3_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_3_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_3_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_3_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_3_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_3_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_3_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_3_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_3_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_3_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_3_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_3_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_3_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_3_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_3_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_3_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_3_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_3_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_3_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_3_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_3_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_3_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_3_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_3_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_3_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_3_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_3_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_3_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_3_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_3_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_3_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_3_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_3_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_3_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_3_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_3_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_3_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_3_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_3_1001 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rst1),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(rst2),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(x1[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(x1[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(x1[11]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(x1[12]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(x1[13]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(x1[14]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(x1[15]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(x1[16]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(x1[17]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(x1[18]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(x1[19]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(x1[1]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(x1[20]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(x1[21]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(x1[22]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(x1[23]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(x1[24]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(x1[25]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(x1[26]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(x1[27]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(x1[28]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(x1[29]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(x1[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(x1[30]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(x1[31]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(x1[3]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(x1[4]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(x1[5]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(x1[6]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(x1[7]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(x1[8]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(x1[9]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(x2[0]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(x2[10]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(x2[11]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(x2[12]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(x2[13]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(x2[14]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(x2[15]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(x2[16]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(x2[17]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(x2[18]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(x2[19]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(x2[1]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(x2[20]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(x2[21]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(x2[22]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(x2[23]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(x2[24]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(x2[25]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(x2[26]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(x2[27]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(x2[28]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(x2[29]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(x2[2]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(x2[30]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(x2[31]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(x2[3]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(x2[4]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(x2[5]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(x2[6]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(x2[7]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(x2[8]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(x2[9]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(y1),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(y2),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 output69 (.A(net69),
    .X(p1));
 sky130_fd_sc_hd__clkbuf_2 output70 (.A(net70),
    .X(p2));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
endmodule
