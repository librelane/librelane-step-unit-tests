../../klayout.streamout/003-success_hybrid/spm.lef