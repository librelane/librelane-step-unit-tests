* NGSPICE file created from aes_core.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__xnor2_2 VGND VPWR Y A B VPB VNB
X0 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_560_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2 VGND B a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X3 Y B a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y a_27_297# a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_474_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X7 VGND A a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X12 a_474_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_560_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VPWR A a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X17 a_560_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__a31o_2 VNB VPB VGND VPWR B1 A1 A2 A3 X
X0 VPWR A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 a_277_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2 a_79_21# B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3 a_277_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_361_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_277_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12675 ps=1.04 w=0.65 l=0.15
X9 a_79_21# A1 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_2 VPWR VGND A X B VPB VNB
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 VGND VPWR VPB VNB CLK D RESET_B Q
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_2 VPB VNB VGND VPWR Y A B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_2 VPWR VGND VPB VNB B2 B1 A1 A2 X
X0 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.102375 ps=0.965 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1575 ps=1.315 w=1 l=0.15
X4 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X5 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X9 a_381_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_2 VGND VPWR VPB VNB S A1 A0 X
X0 VPWR S a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X1 a_591_369# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1312 ps=1.05 w=0.64 l=0.15
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1778 pd=1.415 as=0.135 ps=1.27 w=1 l=0.15
X3 a_79_21# A1 a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1312 pd=1.05 as=0.2288 ps=1.355 w=0.64 l=0.15
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND S a_578_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05775 ps=0.695 w=0.42 l=0.15
X6 a_306_369# a_257_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2288 pd=1.355 as=0.1778 ps=1.415 w=0.64 l=0.15
X7 a_79_21# A0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17325 pd=1.245 as=0.06825 ps=0.745 w=0.42 l=0.15
X8 a_288_47# a_257_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X9 a_257_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_578_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.17325 ps=1.245 w=0.42 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_257_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_2 VNB VPB VGND VPWR X A2 A1 B1 C1
X0 a_79_21# A1 a_348_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.13325 ps=1.06 w=0.65 l=0.15
X1 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.199875 pd=1.265 as=0.091 ps=0.93 w=0.65 l=0.15
X3 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_79_21# C1 a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5 VPWR A2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X6 a_299_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.195 ps=1.39 w=1 l=0.15
X7 a_585_297# B1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_348_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.199875 ps=1.265 w=0.65 l=0.15
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.115375 ps=1.005 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_2 VPWR VGND VPB VNB B D C A X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.91 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_2 Q CLK D VPB VNB VPWR VGND
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X14 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X18 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X19 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X20 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X21 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X22 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2b_2 VPWR VGND VNB VPB A B_N X
X0 VPWR A a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_218_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.15645 ps=1.165 w=0.42 l=0.15
X2 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.15645 pd=1.165 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_300_297# a_27_53# a_218_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 X a_218_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 VPWR a_218_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_218_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X7 VGND a_218_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND A a_218_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_2 VNB VPB VGND VPWR A1 A2 B2 B1 X
X0 a_301_47# B2 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A2 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X2 a_383_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.39 ps=1.78 w=1 l=0.15
X3 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X4 a_301_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X8 VPWR A1 a_579_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X9 a_81_21# B1 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_579_297# A2 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X11 a_81_21# B2 a_383_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 VPB VNB VGND VPWR B Y A
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_2 VPWR VGND VPB VNB C1 B2 B1 A1 A2 X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X1 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1575 ps=1.315 w=1 l=0.15
X3 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.102375 ps=0.965 w=0.65 l=0.15
X6 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X8 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X10 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_2 VPWR VGND X B A VPB VNB
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X6 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X8 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X10 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X11 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X18 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4_2 VNB VPB VGND VPWR D C Y B A
X0 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1 a_471_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=2.84 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_27_47# C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X8 a_277_47# B a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.135 ps=1.27 w=1 l=0.15
X10 Y A a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_277_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X13 a_471_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_2 VGND VPWR VPB VNB B C A X
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4b_2 VNB VPB VGND VPWR A B C Y D_N
X0 VPWR D_N a_694_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_27_297# B a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_474_297# a_694_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_277_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y a_694_21# a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND D_N a_694_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_474_297# C a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y a_694_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_277_297# C a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND a_694_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32ai_2 VPB VNB VGND VPWR A1 A2 Y B1 B2 A3
X0 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X1 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X2 a_475_297# A2 a_729_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3 a_729_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR A1 a_729_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 a_729_297# A2 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_475_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A3 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_2 VNB VPB VGND VPWR A2 A1 Y B1
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_2 VGND VPWR B1 A1 Y A2 VPB VNB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_2 VGND VPWR VNB VPB X C B A_N
X0 a_109_53# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_215_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12715 ps=1.095 w=0.65 l=0.15
X2 a_109_53# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND C a_373_53# VNB sky130_fd_pr__nfet_01v8 ad=0.12715 pd=1.095 as=0.05355 ps=0.675 w=0.42 l=0.15
X4 VGND a_215_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR C a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X6 VPWR a_215_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_215_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X8 a_301_53# a_109_53# a_215_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_215_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_373_53# B a_301_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VPWR a_109_53# a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_2 VPWR VGND VPB VNB X A B
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15575 ps=1.355 w=1 l=0.15
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.355 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111o_2 VNB VPB VGND VPWR A2 A1 B1 C1 X D1
X0 VPWR a_86_235# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND C1 a_86_235# VNB sky130_fd_pr__nfet_01v8 ad=0.121875 pd=1.025 as=0.091 ps=0.93 w=0.65 l=0.15
X2 X a_86_235# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 a_86_235# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.290875 ps=1.545 w=0.65 l=0.15
X4 X a_86_235# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X5 a_715_47# A1 a_86_235# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.108875 ps=0.985 w=0.65 l=0.15
X6 VGND A2 a_715_47# VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 a_499_297# C1 a_427_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X8 VGND a_86_235# X VNB sky130_fd_pr__nfet_01v8 ad=0.290875 pd=1.545 as=0.091 ps=0.93 w=0.65 l=0.15
X9 a_86_235# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.121875 ps=1.025 w=0.65 l=0.15
X10 a_607_297# B1 a_499_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X11 a_427_297# D1 a_86_235# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.41 ps=2.82 w=1 l=0.15
X12 VPWR A1 a_607_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X13 a_607_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_2 VNB VPB VPWR VGND A2 A1 X C1 B1
X0 a_27_47# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3675 pd=1.735 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.23075 pd=2.01 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VPWR A1 a_373_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X4 a_182_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.16535 ps=1.82 w=0.65 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.195 ps=1.39 w=1 l=0.15
X6 a_182_47# B1 a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.16535 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X8 a_373_297# A2 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.3675 ps=1.735 w=1 l=0.15
X9 a_110_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X10 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11 VGND A1 a_182_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_2 VPWR VGND VPB VNB C D_N X A B
X0 a_176_21# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VGND D_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16835 pd=1.495 as=0.135 ps=1.27 w=1 l=0.15
X5 a_555_297# C a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 a_176_21# a_27_53# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1693 ps=1.5 w=1 l=0.15
X8 a_387_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.16835 ps=1.495 w=0.42 l=0.15
X9 a_483_297# B a_387_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 VGND a_27_53# a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 VPWR D_N a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1693 pd=1.5 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.10025 ps=0.985 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311oi_2 VNB VPB VGND VPWR C1 Y B1 A1 A2 A3
X0 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_641_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_297# B1 a_641_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X5 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.17 w=0.65 l=0.15
X11 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X12 a_641_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.0975 ps=0.95 w=0.65 l=0.15
X15 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 Y C1 a_641_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=1.52 w=1 l=0.15
X18 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X19 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_2 VNB VPB VGND VPWR A2 A1 B1 X
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1625 pd=1.15 as=0.1105 ps=0.99 w=0.65 l=0.15
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.1625 ps=1.15 w=0.65 l=0.15
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.1235 ps=1.03 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_2 VGND VPWR VPB VNB X A1 A2 A3 B1
X0 a_108_21# B1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 a_346_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 X a_108_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.26325 ps=2.11 w=0.65 l=0.15
X3 a_108_21# A3 a_430_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_430_297# A2 a_346_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_108_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.175 ps=1.35 w=1 l=0.15
X6 a_346_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND A2 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_108_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.405 ps=2.81 w=1 l=0.15
X9 VPWR B1 a_108_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.2125 ps=1.425 w=1 l=0.15
X10 VGND a_108_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.11375 ps=1 w=0.65 l=0.15
X11 a_346_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_2 B X A C VPWR VGND VPB VNB
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15075 ps=1.345 w=1 l=0.15
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15075 pd=1.345 as=0.074375 ps=0.815 w=0.42 l=0.15
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1304 ps=1.105 w=0.65 l=0.15
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1304 pd=1.105 as=0.05355 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_2 VGND VPWR VPB VNB Y A3 A2 A1 B1
X0 a_281_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1 a_281_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X7 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12675 ps=1.04 w=0.65 l=0.15
X10 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.19825 ps=1.26 w=0.65 l=0.15
X11 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.12675 ps=1.04 w=0.65 l=0.15
X12 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y A3 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.195 ps=1.39 w=1 l=0.15
X15 a_27_297# A2 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311a_2 VPWR VGND VPB VNB X A1 A2 A3 B1 C1
X0 X a_91_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X1 a_91_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X2 a_360_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X3 VPWR B1 a_91_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
X4 a_360_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3125 ps=1.625 w=1 l=0.15
X5 VGND A2 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.11375 ps=1 w=0.65 l=0.15
X6 a_360_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.203125 ps=1.275 w=0.65 l=0.15
X7 VPWR a_91_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND a_91_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 X a_91_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.208 ps=1.94 w=0.65 l=0.15
X10 a_677_47# B1 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X11 a_460_297# A2 a_360_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.175 ps=1.35 w=1 l=0.15
X12 a_91_21# C1 a_677_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X13 a_91_21# A3 a_460_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_2 VNB VPB VGND VPWR C A Y B
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 VPB VNB VPWR VGND Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_2 VNB VPB VGND VPWR B1 B2 A2_N X A1_N
X0 a_294_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.098625 ps=0.98 w=0.42 l=0.15
X1 VPWR A2_N a_295_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2272 pd=1.35 as=0.173 ps=1.4 w=0.64 l=0.15
X2 VPWR B1 a_665_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.18525 ps=1.87 w=0.65 l=0.15
X5 a_581_47# a_295_369# a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X7 a_665_369# B2 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0928 ps=0.93 w=0.64 l=0.15
X8 VGND B2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_295_369# A2_N a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X10 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X11 a_84_21# a_295_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0928 pd=0.93 as=0.2272 ps=1.35 w=0.64 l=0.15
X12 a_295_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.4 as=0.154 ps=1.335 w=0.64 l=0.15
X13 a_581_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_2 VNB VPB VGND VPWR X B1 A2 A1
X0 VPWR A1 a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.16 ps=1.32 w=1 l=0.15
X1 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.4 ps=1.8 w=1 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.089375 ps=0.925 w=0.65 l=0.15
X3 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_470_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.1375 ps=1.275 w=1 l=0.15
X6 a_384_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 a_384_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.104 ps=0.97 w=0.65 l=0.15
X8 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_2 VPB VNB VGND VPWR B1 B2 A2 A1 X C1
X0 VPWR a_38_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A1 a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X2 X a_38_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X3 a_141_47# B2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_497_297# A2 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.3875 ps=1.775 w=1 l=0.15
X5 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR C1 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.325 ps=2.65 w=1 l=0.15
X7 a_237_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1125 pd=1.225 as=0.165 ps=1.33 w=1 l=0.15
X8 a_38_47# B2 a_237_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3875 pd=1.775 as=0.1125 ps=1.225 w=1 l=0.15
X9 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 X a_38_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_141_47# C1 a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.23725 ps=2.03 w=0.65 l=0.15
X12 VGND a_38_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_225_47# B1 a_141_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_2 VPWR VGND VPB VNB C_N X A B
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31oi_2 VNB VPB VPWR VGND B1 Y A1 A2 A3
X0 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.117 ps=1.01 w=0.65 l=0.15
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=1.82 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.175 ps=1.35 w=1 l=0.15
X4 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.41 ps=1.82 w=1 l=0.15
X10 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.18 ps=1.36 w=1 l=0.15
X11 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X13 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0975 ps=0.95 w=0.65 l=0.15
X14 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_2 VNB VPB VGND VPWR B1_N A1 X A2
X0 VPWR A1 a_485_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_485_297# a_297_93# a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 a_297_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.108375 ps=1.01 w=0.42 l=0.15
X3 a_581_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.108375 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_79_21# a_297_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VGND A2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1815 pd=1.51 as=0.14 ps=1.28 w=1 l=0.15
X8 a_297_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1815 ps=1.51 w=0.42 l=0.15
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X10 a_485_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
.ends

.subckt ZI_sky130_fd_sc_hd__nor2_2 VPB VNB VGND VPWR B Y A
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
.ends

.subckt ZI_sky130_fd_sc_hd__a31o_2 VNB VPB VGND VPWR B1 A1 A2 A3 X
X0 VPWR A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 a_277_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2 a_79_21# B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3 a_277_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_361_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_277_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12675 ps=1.04 w=0.65 l=0.15
X9 a_79_21# A1 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__xor2_2 VPWR VGND X B A VPB VNB
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X6 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X8 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X10 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X11 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X18 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__buf_1 VGND VPWR X A VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__dfrtp_2 VGND VPWR VPB VNB CLK D RESET_B Q
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
.ends

.subckt ZI_sky130_fd_sc_hd__or4_2 VPWR VGND VPB VNB B D C A X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.91 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__o21ai_2 VGND VPWR B1 A1 Y A2 VPB VNB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a221o_2 VPWR VGND VPB VNB C1 B2 B1 A1 A2 X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X1 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1575 ps=1.315 w=1 l=0.15
X3 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.102375 ps=0.965 w=0.65 l=0.15
X6 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X8 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X10 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
.ends

.subckt ZI_sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
.ends

.subckt ZI_sky130_fd_sc_hd__xnor2_2 VGND VPWR Y A B VPB VNB
X0 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_560_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2 VGND B a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X3 Y B a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y a_27_297# a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_474_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X7 VGND A a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X12 a_474_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_560_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VPWR A a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X17 a_560_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__or3_2 VGND VPWR VPB VNB B C A X
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a211o_2 VNB VPB VGND VPWR X A2 A1 B1 C1
X0 a_79_21# A1 a_348_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.13325 ps=1.06 w=0.65 l=0.15
X1 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.199875 pd=1.265 as=0.091 ps=0.93 w=0.65 l=0.15
X3 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_79_21# C1 a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5 VPWR A2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X6 a_299_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.195 ps=1.39 w=1 l=0.15
X7 a_585_297# B1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_348_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.199875 ps=1.265 w=0.65 l=0.15
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.115375 ps=1.005 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__o21a_2 VNB VPB VGND VPWR X B1 A2 A1
X0 VPWR A1 a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.16 ps=1.32 w=1 l=0.15
X1 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.4 ps=1.8 w=1 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.089375 ps=0.925 w=0.65 l=0.15
X3 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_470_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.1375 ps=1.275 w=1 l=0.15
X6 a_384_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 a_384_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.104 ps=0.97 w=0.65 l=0.15
X8 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__nor3_2 VPB VNB VGND VPWR A B C Y
X0 Y C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X6 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X10 a_281_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a21oi_2 VNB VPB VGND VPWR A2 A1 Y B1
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__o32a_2 VNB VPB VGND VPWR B1 B2 A3 A2 A1 X
X0 a_429_297# A2 a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND A2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_345_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13975 ps=1.08 w=0.65 l=0.15
X5 a_345_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=1.61 w=1 l=0.15
X6 a_629_297# B2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR B1 a_629_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.19 ps=1.38 w=1 l=0.15
X8 a_79_21# B2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_345_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.1235 ps=1.03 w=0.65 l=0.15
X10 a_79_21# A3 a_429_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_345_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.26 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__and3_2 B X A C VPWR VGND VPB VNB
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15075 ps=1.345 w=1 l=0.15
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15075 pd=1.345 as=0.074375 ps=0.815 w=0.42 l=0.15
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1304 ps=1.105 w=0.65 l=0.15
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1304 pd=1.105 as=0.05355 ps=0.675 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__o211a_2 VNB VPB VPWR VGND A2 A1 X C1 B1
X0 a_27_47# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3675 pd=1.735 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.23075 pd=2.01 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VPWR A1 a_373_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X4 a_182_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.16535 ps=1.82 w=0.65 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.195 ps=1.39 w=1 l=0.15
X6 a_182_47# B1 a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.16535 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X8 a_373_297# A2 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.3675 ps=1.735 w=1 l=0.15
X9 a_110_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X10 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11 VGND A1 a_182_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a21o_2 VNB VPB VGND VPWR A2 A1 B1 X
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1625 pd=1.15 as=0.1105 ps=0.99 w=0.65 l=0.15
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.1625 ps=1.15 w=0.65 l=0.15
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.1235 ps=1.03 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__and2b_2 VNB VPB VPWR VGND A_N X B
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.22895 ps=1.745 w=1 l=0.15
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22895 pd=1.745 as=0.0609 ps=0.71 w=0.42 l=0.15
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__or4b_2 VPWR VGND VPB VNB C D_N X A B
X0 a_176_21# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VGND D_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16835 pd=1.495 as=0.135 ps=1.27 w=1 l=0.15
X5 a_555_297# C a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 a_176_21# a_27_53# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1693 ps=1.5 w=1 l=0.15
X8 a_387_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.16835 ps=1.495 w=0.42 l=0.15
X9 a_483_297# B a_387_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 VGND a_27_53# a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 VPWR D_N a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1693 pd=1.5 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.10025 ps=0.985 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a22o_2 VPWR VGND VPB VNB B2 B1 A1 A2 X
X0 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.102375 ps=0.965 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1575 ps=1.315 w=1 l=0.15
X4 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X5 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X9 a_381_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a2bb2o_2 VNB VPB VGND VPWR B1 B2 A2_N A1_N X
X0 VPWR a_82_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.435 as=0.135 ps=1.27 w=1 l=0.15
X1 a_646_47# B2 a_82_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_574_369# a_313_47# a_82_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0976 pd=0.945 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 a_574_369# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4 VGND a_82_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR B2 a_574_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0976 ps=0.945 w=0.64 l=0.15
X6 X a_82_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 X a_82_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8 a_313_47# A2_N a_313_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.0672 ps=0.85 w=0.64 l=0.15
X9 a_313_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X10 a_313_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.186 ps=1.435 w=0.64 l=0.15
X11 VGND A2_N a_313_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14175 pd=1.095 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_82_21# a_313_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.14175 ps=1.095 w=0.42 l=0.15
X13 VGND B1 a_646_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__o22a_2 VNB VPB VGND VPWR A1 A2 B2 B1 X
X0 a_301_47# B2 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A2 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X2 a_383_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.39 ps=1.78 w=1 l=0.15
X3 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X4 a_301_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X8 VPWR A1 a_579_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X9 a_81_21# B1 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_579_297# A2 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X11 a_81_21# B2 a_383_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__or3b_2 VPWR VGND VPB VNB C_N X A B
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__and2_2 VPWR VGND A X B VPB VNB
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__o41ai_2 VNB VPB VGND VPWR A1 A2 A3 A4 Y B1
X0 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A4 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X4 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_299_297# A3 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X9 a_549_297# A3 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_299_297# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y A4 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_743_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR A1 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_743_297# A2 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_549_297# A2 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X19 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a2111o_2 VNB VPB VGND VPWR A2 A1 B1 C1 X D1
X0 VPWR a_86_235# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND C1 a_86_235# VNB sky130_fd_pr__nfet_01v8 ad=0.121875 pd=1.025 as=0.091 ps=0.93 w=0.65 l=0.15
X2 X a_86_235# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 a_86_235# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.290875 ps=1.545 w=0.65 l=0.15
X4 X a_86_235# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X5 a_715_47# A1 a_86_235# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.108875 ps=0.985 w=0.65 l=0.15
X6 VGND A2 a_715_47# VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 a_499_297# C1 a_427_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X8 VGND a_86_235# X VNB sky130_fd_pr__nfet_01v8 ad=0.290875 pd=1.545 as=0.091 ps=0.93 w=0.65 l=0.15
X9 a_86_235# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.121875 ps=1.025 w=0.65 l=0.15
X10 a_607_297# B1 a_499_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X11 a_427_297# D1 a_86_235# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.41 ps=2.82 w=1 l=0.15
X12 VPWR A1 a_607_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X13 a_607_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__nand2_2 VPB VNB VGND VPWR Y A B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__nand3_2 VNB VPB VGND VPWR C A Y B
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a32o_2 VNB VPB VGND VPWR X A3 A2 B2 B1 A1
X0 VPWR A3 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X2 a_352_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.209625 ps=1.295 w=0.65 l=0.15
X3 a_549_47# A1 a_21_199# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 X a_21_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_21_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.209625 pd=1.295 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13975 ps=1.08 w=0.65 l=0.15
X7 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X8 a_299_297# B1 a_21_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_21_199# B2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND A3 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR a_21_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 X a_21_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_21_199# B1 a_352_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.115375 ps=1.005 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__and3b_2 VGND VPWR VNB VPB X C B A_N
X0 a_109_53# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_215_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12715 ps=1.095 w=0.65 l=0.15
X2 a_109_53# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND C a_373_53# VNB sky130_fd_pr__nfet_01v8 ad=0.12715 pd=1.095 as=0.05355 ps=0.675 w=0.42 l=0.15
X4 VGND a_215_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR C a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X6 VPWR a_215_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_215_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X8 a_301_53# a_109_53# a_215_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_215_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_373_53# B a_301_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VPWR a_109_53# a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__inv_2 VPB VNB VPWR VGND Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__or4bb_2 VPWR VGND VPB VNB B A C_N D_N X
X0 a_398_413# a_206_93# a_316_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1215 pd=1.33 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VPWR a_316_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_316_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X3 X a_316_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X4 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1226 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND a_27_410# a_316_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X7 VGND A a_316_413# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND a_316_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_566_297# B a_494_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05985 pd=0.705 as=0.0441 ps=0.63 w=0.42 l=0.15
X10 a_206_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06195 ps=0.715 w=0.42 l=0.15
X11 a_316_413# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_206_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1226 ps=1.32 w=0.42 l=0.15
X13 a_494_297# a_27_410# a_398_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1215 ps=1.33 w=0.42 l=0.15
X14 a_316_413# a_206_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X15 VPWR A a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.05985 ps=0.705 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__and4b_2 VPWR VGND VNB VPB A_N B C D X
X0 VPWR a_193_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# a_27_413# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.103975 ps=1 w=0.65 l=0.15
X4 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14325 pd=1.33 as=0.06615 ps=0.735 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103975 pd=1 as=0.06195 ps=0.715 w=0.42 l=0.15
X7 VGND a_193_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X8 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X9 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X10 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.14325 ps=1.33 w=1 l=0.15
X11 a_193_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0735 ps=0.77 w=0.42 l=0.15
X13 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__mux2_2 VGND VPWR VPB VNB S A1 A0 X
X0 VPWR S a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X1 a_591_369# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1312 ps=1.05 w=0.64 l=0.15
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1778 pd=1.415 as=0.135 ps=1.27 w=1 l=0.15
X3 a_79_21# A1 a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1312 pd=1.05 as=0.2288 ps=1.355 w=0.64 l=0.15
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND S a_578_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05775 ps=0.695 w=0.42 l=0.15
X6 a_306_369# a_257_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2288 pd=1.355 as=0.1778 ps=1.415 w=0.64 l=0.15
X7 a_79_21# A0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17325 pd=1.245 as=0.06825 ps=0.745 w=0.42 l=0.15
X8 a_288_47# a_257_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X9 a_257_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_578_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.17325 ps=1.245 w=0.42 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_257_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__nand4b_2 VNB VPB VGND VPWR A_N Y B C D
X0 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_465_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND D a_655_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X3 a_215_47# B a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_655_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_655_47# C a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.37 pd=1.74 as=0.135 ps=1.27 w=1 l=0.15
X8 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_465_47# C a_655_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=2.8 as=0.135 ps=1.27 w=1 l=0.15
X13 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.18 ps=1.36 w=1 l=0.15
X14 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.37 ps=1.74 w=1 l=0.15
X17 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__o221a_2 VPB VNB VGND VPWR B1 B2 A2 A1 X C1
X0 VPWR a_38_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A1 a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X2 X a_38_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X3 a_141_47# B2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_497_297# A2 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.3875 ps=1.775 w=1 l=0.15
X5 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR C1 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.325 ps=2.65 w=1 l=0.15
X7 a_237_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1125 pd=1.225 as=0.165 ps=1.33 w=1 l=0.15
X8 a_38_47# B2 a_237_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3875 pd=1.775 as=0.1125 ps=1.225 w=1 l=0.15
X9 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 X a_38_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_141_47# C1 a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.23725 ps=2.03 w=0.65 l=0.15
X12 VGND a_38_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_225_47# B1 a_141_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__and4_2 VNB VPB VGND VPWR X D C B A
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.27995 ps=1.615 w=1 l=0.15
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.06195 ps=0.715 w=0.42 l=0.15
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.17515 ps=1.265 w=0.65 l=0.15
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.07455 ps=0.775 w=0.42 l=0.15
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a41oi_2 VNB VPB VPWR VGND A4 A3 A2 A1 B1 Y
X0 a_149_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_757_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_757_47# A3 a_567_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR A3 a_149_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=1.77 as=0.145 ps=1.29 w=1 l=0.15
X4 Y B1 a_149_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_567_47# A3 a_757_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VGND A4 a_757_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A4 a_149_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_149_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_317_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_317_47# A2 a_567_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_149_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.385 ps=1.77 w=1 l=0.15
X13 a_149_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A1 a_317_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 VPWR A2 a_149_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_567_47# A2 a_317_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_149_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VPWR A1 a_149_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__or2b_2 VPWR VGND VNB VPB A B_N X
X0 VPWR A a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_218_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.15645 ps=1.165 w=0.42 l=0.15
X2 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.15645 pd=1.165 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_300_297# a_27_53# a_218_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 X a_218_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 VPWR a_218_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_218_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X7 VGND a_218_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND A a_218_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__or2_2 VPWR VGND VPB VNB X A B
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15575 ps=1.355 w=1 l=0.15
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.355 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__o22ai_2 VPB VNB VGND VPWR A1 A2 Y B2 B1
X0 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_475_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR A1 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.26975 pd=1.48 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12 a_475_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 Y A2 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X14 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.26975 ps=1.48 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a41o_2 VNB VPB VGND VPWR X A1 A2 A3 A4 B1
X0 a_381_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A2 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X2 a_465_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_549_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13975 ps=1.08 w=0.65 l=0.15
X7 a_381_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A4 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_381_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 a_79_21# A1 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__o2bb2a_2 VNB VPB VGND VPWR B1 B2 A2_N X A1_N
X0 a_294_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.098625 ps=0.98 w=0.42 l=0.15
X1 VPWR A2_N a_295_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2272 pd=1.35 as=0.173 ps=1.4 w=0.64 l=0.15
X2 VPWR B1 a_665_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.18525 ps=1.87 w=0.65 l=0.15
X5 a_581_47# a_295_369# a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X7 a_665_369# B2 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0928 ps=0.93 w=0.64 l=0.15
X8 VGND B2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_295_369# A2_N a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X10 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X11 a_84_21# a_295_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0928 pd=0.93 as=0.2272 ps=1.35 w=0.64 l=0.15
X12 a_295_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.4 as=0.154 ps=1.335 w=0.64 l=0.15
X13 a_581_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__o41a_2 VNB VPB VGND VPWR A1 A2 A3 A4 B1 X
X0 VGND A2 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.11375 ps=1 w=0.65 l=0.15
X1 a_496_297# A4 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.3025 ps=1.605 w=1 l=0.15
X2 a_393_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.115375 ps=1.005 w=0.65 l=0.15
X3 VPWR A1 a_697_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=2.82 as=0.175 ps=1.35 w=1 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3025 pd=1.605 as=0.305 ps=1.61 w=1 l=0.15
X7 VGND A4 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.118625 ps=1.015 w=0.65 l=0.15
X8 a_697_297# A2 a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X9 a_393_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2665 pd=2.12 as=0.11375 ps=1 w=0.65 l=0.15
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_393_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.208 ps=1.94 w=0.65 l=0.15
X12 a_597_297# A3 a_496_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.1775 ps=1.355 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__o211ai_2 VNB VPB VGND VPWR Y B1 A2 A1 C1
X0 a_286_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2 a_286_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X3 Y A2 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 VGND A1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X6 VGND A2 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 a_487_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_27_47# B1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR A1 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X13 a_487_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14 a_286_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__o31ai_2 VGND VPWR VPB VNB Y A3 A2 A1 B1
X0 a_281_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1 a_281_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X7 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12675 ps=1.04 w=0.65 l=0.15
X10 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.19825 ps=1.26 w=0.65 l=0.15
X11 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.12675 ps=1.04 w=0.65 l=0.15
X12 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y A3 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.195 ps=1.39 w=1 l=0.15
X15 a_27_297# A2 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__o31a_2 VGND VPWR VPB VNB X A1 A2 A3 B1
X0 a_108_21# B1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 a_346_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 X a_108_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.26325 ps=2.11 w=0.65 l=0.15
X3 a_108_21# A3 a_430_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_430_297# A2 a_346_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_108_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.175 ps=1.35 w=1 l=0.15
X6 a_346_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND A2 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_108_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.405 ps=2.81 w=1 l=0.15
X9 VPWR B1 a_108_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.2125 ps=1.425 w=1 l=0.15
X10 VGND a_108_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.11375 ps=1 w=0.65 l=0.15
X11 a_346_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a311o_2 VPB VNB VGND VPWR C1 B1 A1 A2 A3 X
X0 a_79_21# C1 a_635_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.21 ps=1.42 w=1 l=0.15
X1 VPWR A2 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.17 ps=1.34 w=1 l=0.15
X2 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.13325 ps=1.06 w=0.65 l=0.15
X3 a_417_47# A2 a_319_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.1105 ps=0.99 w=0.65 l=0.15
X4 a_79_21# A1 a_417_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12025 ps=1.02 w=0.65 l=0.15
X5 a_319_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.156 ps=1.13 w=0.65 l=0.15
X6 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.24 pd=1.48 as=0.135 ps=1.27 w=1 l=0.15
X7 a_319_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.185 ps=1.37 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.156 pd=1.13 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_319_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.34 as=0.24 ps=1.48 w=1 l=0.15
X10 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13975 ps=1.08 w=0.65 l=0.15
X11 a_635_297# B1 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.21 ps=1.42 w=1 l=0.15
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__nand3b_2 VNB VPB VGND VPWR A_N C B Y
X0 a_408_47# B a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_408_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y a_27_47# a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17575 pd=1.395 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND C a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 a_218_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11975 ps=1.045 w=0.65 l=0.15
X7 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_218_47# B a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.17575 ps=1.395 w=1 l=0.15
X12 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11975 pd=1.045 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__nor3b_2 VPB VNB VGND VPWR A Y C_N B
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND a_531_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR C_N a_531_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9 a_281_297# a_531_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X10 Y a_531_21# a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 VGND C_N a_531_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X13 Y a_531_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a22oi_2 VPWR VGND VPB VNB B2 B1 Y A1 A2
X0 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_467_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_467_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_109_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__o311a_2 VPWR VGND VPB VNB X A1 A2 A3 B1 C1
X0 X a_91_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X1 a_91_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X2 a_360_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X3 VPWR B1 a_91_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
X4 a_360_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3125 ps=1.625 w=1 l=0.15
X5 VGND A2 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.11375 ps=1 w=0.65 l=0.15
X6 a_360_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.203125 ps=1.275 w=0.65 l=0.15
X7 VPWR a_91_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND a_91_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 X a_91_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.208 ps=1.94 w=0.65 l=0.15
X10 a_677_47# B1 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X11 a_460_297# A2 a_360_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.175 ps=1.35 w=1 l=0.15
X12 a_91_21# C1 a_677_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X13 a_91_21# A3 a_460_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a31oi_2 VNB VPB VPWR VGND B1 Y A1 A2 A3
X0 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.117 ps=1.01 w=0.65 l=0.15
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=1.82 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.175 ps=1.35 w=1 l=0.15
X4 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.41 ps=1.82 w=1 l=0.15
X10 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.18 ps=1.36 w=1 l=0.15
X11 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X13 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0975 ps=0.95 w=0.65 l=0.15
X14 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__and4bb_2 VNB VPB VGND VPWR A_N X C D B_N
X0 a_174_21# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1 a_174_21# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.33075 ps=1.705 w=0.42 l=0.15
X2 a_476_47# a_27_47# a_174_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33075 pd=1.705 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X5 a_548_47# a_505_280# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8 VPWR D a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND D a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 VPWR a_505_280# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X11 a_505_280# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X12 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_505_280# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X14 a_639_47# C a_548_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X15 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__dfstp_2 VPB VNB VPWR VGND Q SET_B D CLK
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.06705 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_1136_413# a_193_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X3 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06705 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X5 a_1228_47# a_27_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X6 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X8 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12495 pd=1.175 as=0.2184 ps=2.2 w=0.84 l=0.15
X10 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X11 VPWR a_1602_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1028_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VGND a_1602_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_1028_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.12495 ps=1.175 w=0.42 l=0.15
X18 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1028_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X20 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X21 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_1028_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0441 ps=0.63 w=0.42 l=0.15
X23 VPWR a_1178_261# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X24 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 a_1178_261# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2226 pd=2.21 as=0.12075 ps=1.165 w=0.84 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_1300_47# a_1178_261# a_1228_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X28 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X29 a_1178_261# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1404 pd=1.6 as=0.1137 ps=1.01 w=0.54 l=0.15
X30 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X31 VPWR SET_B a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12075 pd=1.165 as=0.1092 ps=1.36 w=0.42 l=0.15
X32 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X33 VGND SET_B a_1300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1137 pd=1.01 as=0.0441 ps=0.63 w=0.42 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a221oi_2 VNB VPB VGND VPWR A2 A1 B1 B2 Y C1
X0 Y B1 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_301_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_301_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND B2 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A1 a_735_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_297# B2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR A1 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_735_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_301_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1755 ps=1.84 w=0.65 l=0.15
X12 VPWR A2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X13 a_383_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X14 a_383_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_735_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X16 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X17 a_301_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X18 a_735_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B1 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__o2111a_2 VPB VNB VGND VPWR X D1 C1 B1 A2 A1
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 a_80_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.365 ps=1.73 w=1 l=0.15
X3 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VPWR C1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.14 ps=1.28 w=1 l=0.15
X5 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X6 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X7 a_674_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X8 a_386_47# D1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X9 VPWR A1 a_674_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.195 ps=1.39 w=1 l=0.15
X10 a_566_47# B1 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X11 VGND A2 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X12 a_566_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X13 a_458_47# C1 a_386_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a21bo_2 VNB VPB VGND VPWR B1_N A1 X A2
X0 VPWR A1 a_485_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_485_297# a_297_93# a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 a_297_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.108375 ps=1.01 w=0.42 l=0.15
X3 a_581_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.108375 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_79_21# a_297_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VGND A2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1815 pd=1.51 as=0.14 ps=1.28 w=1 l=0.15
X8 a_297_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1815 ps=1.51 w=0.42 l=0.15
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X10 a_485_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__o221ai_2 VNB VPB VGND VPWR Y B1 B2 A2 A1 C1
X0 Y A2 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_300_47# B2 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 a_300_47# B1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_300_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_734_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X7 a_28_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y C1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR B1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X11 a_382_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_28_47# B1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_28_47# B2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X15 Y B2 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VPWR A1 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND A2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_382_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X19 a_734_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a32oi_2 VNB VPB VGND VPWR B2 B1 Y A1 A2 A3
X0 Y A1 a_478_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.3775 ps=1.755 w=1 l=0.15
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.305 ps=1.61 w=1 l=0.15
X3 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.335 ps=1.67 w=1 l=0.15
X4 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.1375 ps=1.275 w=1 l=0.15
X5 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3775 pd=1.755 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_478_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_478_47# A2 a_730_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND A3 a_730_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12025 ps=1.02 w=0.65 l=0.15
X10 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_730_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.20475 ps=1.93 w=0.65 l=0.15
X16 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.15 ps=1.3 w=1 l=0.15
X18 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X19 a_730_47# A2 a_478_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__nand4_2 VNB VPB VGND VPWR D C Y B A
X0 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1 a_471_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=2.84 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_27_47# C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X8 a_277_47# B a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.135 ps=1.27 w=1 l=0.15
X10 Y A a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_277_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X13 a_471_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a211oi_2 VPWR VGND VPB VNB A2 A1 Y B1 C1
X0 VGND A2 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR A1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_37_297# B1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_485_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_292_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VPWR A2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_485_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X11 a_37_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 Y A1 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X13 Y C1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14 a_292_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15 a_292_297# B1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__a2111oi_2 VNB VPB VGND VPWR A1 A2 D1 C1 B1 Y
X0 a_467_297# B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X1 a_287_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR A2 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X3 a_923_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.112125 ps=0.995 w=0.65 l=0.15
X4 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X5 a_28_297# B1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X7 a_28_297# C1 a_287_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X8 Y A1 a_923_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND A2 a_684_47# VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17875 ps=1.2 w=0.65 l=0.15
X10 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.105625 ps=0.975 w=0.65 l=0.15
X12 Y D1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_467_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=2.67 as=0.16 ps=1.32 w=1 l=0.15
X14 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.12675 ps=1.04 w=0.65 l=0.15
X16 VPWR A1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X17 a_115_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X18 a_467_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 a_684_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.2 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt ZI_sky130_fd_sc_hd__nor4_2 VNB VPB VGND VPWR B D Y A C
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_475_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y D a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12 a_475_297# C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_281_297# C a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X14 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X15 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
.ends

.subckt aes_decipher_block block[0] block[100] block[101] block[102] block[103] block[104]
+ block[105] block[106] block[107] block[108] block[109] block[10] block[110] block[111]
+ block[112] block[113] block[114] block[115] block[116] block[117] block[118] block[119]
+ block[11] block[120] block[121] block[122] block[123] block[124] block[125] block[126]
+ block[127] block[12] block[13] block[14] block[15] block[16] block[17] block[18]
+ block[19] block[1] block[20] block[21] block[22] block[23] block[24] block[25] block[26]
+ block[27] block[28] block[29] block[2] block[30] block[31] block[32] block[33] block[34]
+ block[35] block[36] block[37] block[38] block[39] block[3] block[40] block[41] block[42]
+ block[43] block[44] block[45] block[46] block[47] block[48] block[49] block[4] block[50]
+ block[51] block[52] block[53] block[54] block[55] block[56] block[57] block[58]
+ block[59] block[5] block[60] block[61] block[62] block[63] block[64] block[65] block[66]
+ block[67] block[68] block[69] block[6] block[70] block[71] block[72] block[73] block[74]
+ block[75] block[76] block[77] block[78] block[79] block[7] block[80] block[81] block[82]
+ block[83] block[84] block[85] block[86] block[87] block[88] block[89] block[8] block[90]
+ block[91] block[92] block[93] block[94] block[95] block[96] block[97] block[98]
+ block[99] block[9] clk keylen new_block[0] new_block[100] new_block[101] new_block[102]
+ new_block[103] new_block[104] new_block[105] new_block[106] new_block[107] new_block[108]
+ new_block[109] new_block[10] new_block[110] new_block[111] new_block[112] new_block[113]
+ new_block[114] new_block[115] new_block[116] new_block[117] new_block[118] new_block[119]
+ new_block[11] new_block[120] new_block[121] new_block[122] new_block[123] new_block[124]
+ new_block[125] new_block[126] new_block[127] new_block[12] new_block[13] new_block[14]
+ new_block[15] new_block[16] new_block[17] new_block[18] new_block[19] new_block[1]
+ new_block[20] new_block[21] new_block[22] new_block[23] new_block[24] new_block[25]
+ new_block[26] new_block[27] new_block[28] new_block[29] new_block[2] new_block[30]
+ new_block[31] new_block[32] new_block[33] new_block[34] new_block[35] new_block[36]
+ new_block[37] new_block[38] new_block[39] new_block[3] new_block[40] new_block[41]
+ new_block[42] new_block[43] new_block[44] new_block[45] new_block[46] new_block[47]
+ new_block[48] new_block[49] new_block[4] new_block[50] new_block[51] new_block[52]
+ new_block[53] new_block[54] new_block[55] new_block[56] new_block[57] new_block[58]
+ new_block[59] new_block[5] new_block[60] new_block[61] new_block[62] new_block[63]
+ new_block[64] new_block[65] new_block[66] new_block[67] new_block[68] new_block[69]
+ new_block[6] new_block[70] new_block[71] new_block[72] new_block[73] new_block[74]
+ new_block[75] new_block[76] new_block[77] new_block[78] new_block[79] new_block[7]
+ new_block[80] new_block[81] new_block[82] new_block[83] new_block[84] new_block[85]
+ new_block[86] new_block[87] new_block[88] new_block[89] new_block[8] new_block[90]
+ new_block[91] new_block[92] new_block[93] new_block[94] new_block[95] new_block[96]
+ new_block[97] new_block[98] new_block[99] new_block[9] next ready reset_n round[0]
+ round[1] round[2] round[3] round_key[0] round_key[100] round_key[101] round_key[102]
+ round_key[103] round_key[104] round_key[105] round_key[106] round_key[107] round_key[108]
+ round_key[109] round_key[10] round_key[110] round_key[111] round_key[112] round_key[113]
+ round_key[114] round_key[115] round_key[116] round_key[117] round_key[118] round_key[119]
+ round_key[11] round_key[120] round_key[121] round_key[122] round_key[123] round_key[124]
+ round_key[125] round_key[126] round_key[127] round_key[12] round_key[13] round_key[14]
+ round_key[15] round_key[16] round_key[17] round_key[18] round_key[19] round_key[1]
+ round_key[20] round_key[21] round_key[22] round_key[23] round_key[24] round_key[25]
+ round_key[26] round_key[27] round_key[28] round_key[29] round_key[2] round_key[30]
+ round_key[31] round_key[32] round_key[33] round_key[34] round_key[35] round_key[36]
+ round_key[37] round_key[38] round_key[39] round_key[3] round_key[40] round_key[41]
+ round_key[42] round_key[43] round_key[44] round_key[45] round_key[46] round_key[47]
+ round_key[48] round_key[49] round_key[4] round_key[50] round_key[51] round_key[52]
+ round_key[53] round_key[54] round_key[55] round_key[56] round_key[57] round_key[58]
+ round_key[59] round_key[5] round_key[60] round_key[61] round_key[62] round_key[63]
+ round_key[64] round_key[65] round_key[66] round_key[67] round_key[68] round_key[69]
+ round_key[6] round_key[70] round_key[71] round_key[72] round_key[73] round_key[74]
+ round_key[75] round_key[76] round_key[77] round_key[78] round_key[79] round_key[7]
+ round_key[80] round_key[81] round_key[82] round_key[83] round_key[84] round_key[85]
+ round_key[86] round_key[87] round_key[88] round_key[89] round_key[8] round_key[90]
+ round_key[91] round_key[92] round_key[93] round_key[94] round_key[95] round_key[96]
+ round_key[97] round_key[98] round_key[99] round_key[9] VPWR VGND
XFILLER_0_94_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7963_ VPWR VGND VGND VPWR _0808_ _3356_ _4090_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_96_409 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6914_ VGND VPWR VGND VPWR _2185_ _2339_ _2233_ _2297_ _2367_ ZI_sky130_fd_sc_hd__a31o_2
X_7894_ VPWR VGND _3293_ block[111] round_key[111] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6845_ VGND VPWR _2299_ _2141_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6776_ VGND VPWR _2230_ _2213_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_76_188 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_9_499 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5727_ VPWR VGND _1192_ _0907_ _0795_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8515_ VGND VPWR VPWR VGND clk _0117_ reset_n new_block[10] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_91_169 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8446_ VGND VPWR VPWR VGND clk _0048_ reset_n new_block[69] ZI_sky130_fd_sc_hd__dfrtp_2
X_5658_ VPWR VGND VPWR VGND _1106_ _1123_ _1110_ _0824_ _1124_ ZI_sky130_fd_sc_hd__or4_2
X_5589_ VGND VPWR _4103_ _4090_ _1056_ _1055_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
X_8377_ VPWR VGND VPWR VGND _3521_ _4093_ _3729_ _0169_ _1574_ _3730_ ZI_sky130_fd_sc_hd__a221o_2
X_4609_ VPWR VGND VGND VPWR _4145_ _4146_ _4008_ ZI_sky130_fd_sc_hd__nor2_2
X_7328_ VPWR VGND VPWR VGND _2757_ _2774_ _2763_ _2746_ _2775_ ZI_sky130_fd_sc_hd__or4_2
X_7259_ VPWR VGND VPWR VGND _2383_ _2706_ _2568_ _2332_ _2707_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_99_214 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_99_225 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_68_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_68_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_67_188 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_23_203 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_51_523 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_23_269 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_3_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4960_ VGND VPWR _0433_ _0430_ _0432_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_133 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4891_ VPWR VGND VGND VPWR _4083_ _0365_ _4082_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_13_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_104_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6630_ VGND VPWR VPWR VGND _2078_ _2083_ _3775_ _2084_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_73_125 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6561_ VGND VPWR VGND VPWR _2016_ _1546_ _1375_ _1867_ _2015_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_13_62 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_73_169 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8300_ VGND VPWR _3660_ _0802_ _1139_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5512_ VGND VPWR VGND VPWR _0980_ _0841_ _0825_ _0975_ ZI_sky130_fd_sc_hd__o21a_2
X_6492_ VPWR VGND _1949_ _1762_ _1574_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5443_ VPWR VGND _0912_ round_key[54] new_block[54] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8231_ VGND VPWR _3598_ _0383_ _0477_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5374_ VPWR VGND VPWR VGND _0761_ _0644_ _0765_ _0618_ _0634_ _0843_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_112_477 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8162_ VGND VPWR _3536_ _0296_ _0307_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7113_ VPWR VGND _2564_ block[123] round_key[123] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4325_ VPWR VGND VGND VPWR _3832_ _3835_ _3836_ _3863_ ZI_sky130_fd_sc_hd__nor3_2
X_8093_ VPWR VGND _3473_ _2776_ _2416_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7044_ VPWR VGND _2496_ block[122] round_key[122] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4256_ VPWR VGND VGND VPWR _3793_ _3794_ _3787_ ZI_sky130_fd_sc_hd__nor2_2
X_7946_ VGND VPWR VGND VPWR _3338_ _3332_ _3340_ _3339_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_77_442 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7877_ VGND VPWR VGND VPWR _3240_ new_block[45] _3277_ _3275_ _1181_ _0088_ ZI_sky130_fd_sc_hd__o32a_2
X_6828_ VGND VPWR _2282_ _2281_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_45_350 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6759_ VGND VPWR _2213_ _2212_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_33_556 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_45_383 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8429_ VGND VPWR VPWR VGND clk _0031_ reset_n new_block[116] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_228 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_18_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_50_16 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_36_372 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_51_397 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_59_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5090_ sword_ctr_reg\[1\] _0560_ sword_ctr_reg\[0\] new_block[14] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
X_5992_ VGND VPWR VGND VPWR _1454_ _1453_ _1426_ _1340_ ZI_sky130_fd_sc_hd__o21a_2
X_7800_ VGND VPWR VPWR VGND _3206_ _3201_ _3208_ _3118_ _3207_ ZI_sky130_fd_sc_hd__o211a_2
X_7731_ VGND VPWR _3145_ _1683_ _3144_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4943_ VPWR VGND VPWR VGND _4048_ _0415_ _0412_ _4024_ _0416_ ZI_sky130_fd_sc_hd__or4_2
X_7662_ VGND VPWR VGND VPWR _3079_ _0444_ _3081_ _3082_ ZI_sky130_fd_sc_hd__a21o_2
X_6613_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] _2067_ new_block[95] ZI_sky130_fd_sc_hd__and2b_2
X_4874_ VPWR VGND VPWR VGND _0346_ _0347_ _0348_ _0344_ _0345_ ZI_sky130_fd_sc_hd__or4b_2
XFILLER_0_6_222 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_62_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7593_ VGND VPWR VGND VPWR _3016_ _0444_ _3018_ _3019_ ZI_sky130_fd_sc_hd__a21o_2
XPHY_EDGE_ROW_104_Left_217 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6544_ VPWR VGND _2000_ _1819_ _1762_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_61_128 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6475_ _1390_ _1932_ _1335_ _1332_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5426_ VPWR VGND VPWR VGND _0607_ _0763_ _0601_ _0748_ _0895_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_71_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8214_ VGND VPWR _3583_ _0168_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_100_414 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5357_ _0734_ _0826_ _0654_ _0771_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8145_ VGND VPWR _3521_ _3458_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5288_ VGND VPWR VPWR VGND _0757_ _0628_ _0758_ _0580_ _0630_ ZI_sky130_fd_sc_hd__o211a_2
X_8076_ VGND VPWR VGND VPWR _4099_ _3777_ _0001_ _3751_ _3458_ ZI_sky130_fd_sc_hd__a2bb2o_2
X_4308_ VGND VPWR VPWR VGND _3827_ _3829_ _3832_ _3846_ ZI_sky130_fd_sc_hd__or3_2
X_7027_ VGND VPWR VGND VPWR _2479_ _2194_ _2196_ _2478_ _2198_ ZI_sky130_fd_sc_hd__a211o_2
X_4239_ VGND VPWR _0007_ _3780_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_69_217 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7929_ VGND VPWR _3324_ _3320_ _3323_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_514 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_92_242 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_37_169 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_108_569 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_29_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_103_296 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_45_16 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_44_607 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_71_404 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_9_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Right_104 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4590_ VGND VPWR VGND VPWR _3905_ _4125_ _3993_ _4035_ _4127_ ZI_sky130_fd_sc_hd__o22a_2
XFILLER_0_3_225 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_10_74 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_10_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6260_ VGND VPWR _1719_ _1655_ _1720_ _1447_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
X_6191_ VPWR VGND VPWR VGND _1414_ _1652_ _1352_ _1362_ ZI_sky130_fd_sc_hd__or3b_2
X_5211_ VGND VPWR VPWR VGND _0660_ _0680_ _0647_ _0681_ ZI_sky130_fd_sc_hd__or3_2
X_5142_ VPWR VGND _0531_ _0612_ _0600_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5073_ VGND VPWR VGND VPWR _0538_ _0539_ _0540_ _0541_ _0543_ _0542_ ZI_sky130_fd_sc_hd__o41ai_2
XFILLER_0_35_93 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5975_ VPWR VGND VGND VPWR _1436_ _1437_ _1388_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_19_125 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7714_ VPWR VGND _3130_ block[94] round_key[94] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4926_ VGND VPWR VGND VPWR _4010_ _3869_ _3931_ _0399_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_7_531 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_19_169 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4857_ VGND VPWR VGND VPWR _3954_ _3872_ _4052_ _4141_ _0331_ ZI_sky130_fd_sc_hd__o22a_2
X_7645_ VGND VPWR _3066_ _0155_ _3065_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7576_ VGND VPWR _3003_ _3001_ _3002_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_517 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6527_ VGND VPWR VPWR VGND _1936_ _1982_ _1977_ _1983_ ZI_sky130_fd_sc_hd__or3_2
X_4788_ VPWR VGND VPWR VGND _3985_ _0262_ _4044_ _4138_ _0263_ ZI_sky130_fd_sc_hd__or4_2
X_6458_ VGND VPWR VGND VPWR _1616_ _1527_ _1483_ _1478_ _1915_ _1467_ ZI_sky130_fd_sc_hd__a2111o_2
X_6389_ VGND VPWR VGND VPWR _1549_ _1609_ _1847_ _1371_ ZI_sky130_fd_sc_hd__a21oi_2
X_5409_ VGND VPWR VGND VPWR _0877_ _0577_ _0579_ _0606_ _0878_ ZI_sky130_fd_sc_hd__a31o_2
X_8128_ VPWR VGND _3505_ _3026_ _0363_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8059_ VGND VPWR VGND VPWR _3152_ new_block[62] _3442_ _3435_ _2731_ _0105_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_85_518 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_38_489 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_56_37 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_56_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5760_ VPWR VGND VPWR VGND _1220_ _1223_ _1222_ _1218_ _1224_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_17_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4711_ VGND VPWR VGND VPWR _4154_ _0186_ _0187_ _4046_ ZI_sky130_fd_sc_hd__a21oi_2
X_5691_ VPWR VGND VPWR VGND _1027_ _1155_ _1153_ _1150_ _1156_ ZI_sky130_fd_sc_hd__or4_2
X_7430_ VPWR VGND VGND VPWR _2869_ _2870_ _0158_ ZI_sky130_fd_sc_hd__nor2_2
X_4642_ VGND VPWR VGND VPWR _3933_ _4016_ _3999_ _4178_ _4179_ ZI_sky130_fd_sc_hd__o22a_2
XFILLER_0_112_53 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_21_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_25_651 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7361_ VPWR VGND VGND VPWR _2806_ _0797_ _2805_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_24_172 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_112_97 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4573_ VGND VPWR _4110_ _4109_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_4_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6312_ VGND VPWR VGND VPWR _1009_ new_block[114] _1771_ _1768_ _1750_ _0029_ ZI_sky130_fd_sc_hd__o32a_2
X_7292_ VPWR VGND _2740_ _2739_ _2738_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6243_ VPWR VGND VPWR VGND _1449_ _1702_ _1699_ _1387_ _1703_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_97_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6174_ VPWR VGND _1394_ _1635_ _1426_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5125_ _0593_ _0595_ _3914_ _0594_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5056_ VGND VPWR VGND VPWR new_block[9] sword_ctr_reg\[0\] _0526_ sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__nand3_2
X_5958_ _1295_ _1420_ _1400_ _1381_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_62_91 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4909_ VPWR VGND _0383_ _0382_ _4061_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5889_ VGND VPWR _1351_ _1350_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7628_ VPWR VGND _3051_ block[119] round_key[119] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7559_ VGND VPWR _2987_ _2639_ _2687_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_153 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_30_197 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_101_586 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_26_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_97_131 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_97_142 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_58_507 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_58_529 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_53_201 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_108_141 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_109_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_53_234 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_81_554 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_13_109 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_34_492 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_83_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_89_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6930_ VGND VPWR VGND VPWR _2383_ _2213_ _2339_ _2345_ _2228_ _2382_ ZI_sky130_fd_sc_hd__a32o_2
X_6861_ VPWR VGND _2315_ _1241_ _1198_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_107_86 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5812_ VGND VPWR _1275_ _1271_ _1274_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_604 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6792_ VGND VPWR _2246_ _2245_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5743_ VGND VPWR VPWR VGND _1205_ _1206_ _1120_ _1207_ ZI_sky130_fd_sc_hd__or3_2
X_8531_ VGND VPWR VPWR VGND clk _0133_ reset_n new_block[26] ZI_sky130_fd_sc_hd__dfrtp_2
X_5674_ VGND VPWR _1140_ _1137_ _1139_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8462_ VGND VPWR VPWR VGND clk _0064_ reset_n new_block[85] ZI_sky130_fd_sc_hd__dfrtp_2
X_7413_ VPWR VGND VGND VPWR _2854_ _2847_ _2853_ ZI_sky130_fd_sc_hd__nand2_2
X_4625_ VPWR VGND VPWR VGND _4018_ _4161_ _4158_ _4011_ _4162_ ZI_sky130_fd_sc_hd__or4_2
X_8393_ VPWR VGND VGND VPWR _3744_ _3742_ _3743_ ZI_sky130_fd_sc_hd__nand2_2
X_7344_ VPWR VGND _2790_ _0810_ _0794_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4556_ VGND VPWR _4094_ _4093_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_4_386 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_13_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_12_197 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4487_ VPWR VGND VGND VPWR _4025_ _3881_ _3959_ ZI_sky130_fd_sc_hd__nand2_2
X_7275_ VPWR VGND VPWR VGND _2609_ _2177_ _2235_ _2096_ _2141_ _2723_ ZI_sky130_fd_sc_hd__a221o_2
X_6226_ VGND VPWR _1687_ _1678_ _1686_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6157_ VGND VPWR VGND VPWR _1617_ _1515_ _1474_ _1616_ _1618_ ZI_sky130_fd_sc_hd__a31o_2
X_5108_ VGND VPWR VGND VPWR _0543_ _0537_ _3850_ _0578_ ZI_sky130_fd_sc_hd__a21o_2
X_6088_ VPWR VGND VGND VPWR _1549_ _1550_ _1547_ ZI_sky130_fd_sc_hd__nor2_2
X_5039_ VGND VPWR VGND VPWR _3896_ _3933_ _0510_ _3870_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_94_134 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_67_337 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_94_178 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_106_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_106_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_37_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_53_16 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_86_602 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_86_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_189 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_41_204 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4410_ VGND VPWR _3948_ _3857_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5390_ VGND VPWR _0859_ _0741_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_41_259 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_111_169 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4341_ VGND VPWR _3879_ _3773_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_10_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7060_ VGND VPWR VGND VPWR _2510_ _2219_ _2199_ _2178_ _2511_ ZI_sky130_fd_sc_hd__a31o_2
X_4272_ VGND VPWR VGND VPWR _3810_ sword_ctr_reg\[0\] new_block[67] sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__and3b_2
X_6011_ VGND VPWR _1473_ _1472_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7962_ VPWR VGND _3355_ block[85] round_key[85] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6913_ VGND VPWR VPWR VGND _2359_ _2365_ _2357_ _2366_ ZI_sky130_fd_sc_hd__or3_2
X_7893_ VPWR VGND VPWR VGND _3292_ _0799_ ZI_sky130_fd_sc_hd__inv_2
XFILLER_0_49_337 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6844_ VGND VPWR VGND VPWR _2298_ _2297_ _2282_ _2178_ ZI_sky130_fd_sc_hd__o21a_2
X_6775_ VGND VPWR _2229_ _2228_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_92_638 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5726_ VGND VPWR _1191_ _1183_ _1190_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8514_ VGND VPWR VPWR VGND clk _0116_ reset_n new_block[9] ZI_sky130_fd_sc_hd__dfrtp_2
X_8445_ VGND VPWR VPWR VGND clk _0047_ reset_n new_block[68] ZI_sky130_fd_sc_hd__dfrtp_2
X_5657_ VPWR VGND VPWR VGND _1115_ _1122_ _1119_ _0743_ _1123_ ZI_sky130_fd_sc_hd__or4_2
X_5588_ VGND VPWR _1055_ round_key[107] new_block[107] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_114 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8376_ VPWR VGND _3729_ block[29] round_key[29] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4608_ VGND VPWR VGND VPWR _4115_ _4141_ _3955_ _4052_ _4145_ ZI_sky130_fd_sc_hd__o22a_2
X_7327_ VPWR VGND VPWR VGND _2659_ _2773_ _2765_ _2764_ _2774_ ZI_sky130_fd_sc_hd__or4_2
X_4539_ VPWR VGND _4077_ round_key[72] new_block[72] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7258_ VPWR VGND VPWR VGND _2665_ _2194_ _2246_ _2097_ _2150_ _2706_ ZI_sky130_fd_sc_hd__a221o_2
X_6209_ VGND VPWR VGND VPWR _1462_ _1609_ _1670_ _1371_ ZI_sky130_fd_sc_hd__a21oi_2
X_7189_ VGND VPWR _2639_ _1006_ _1280_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_68_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_68_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_23_215 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_23_237 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_48_16 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_59_613 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_86_421 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_59_646 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4890_ VGND VPWR _4103_ _4090_ _0364_ _0363_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_17_Left_130 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6560_ VGND VPWR VGND VPWR _2015_ _1456_ _1419_ _1361_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_27_532 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_104_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_73_159 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5511_ _0688_ _0979_ _0630_ _0699_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6491_ VGND VPWR _1948_ _1757_ _1947_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5442_ VPWR VGND _0911_ round_key[49] new_block[49] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_112_434 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8230_ VGND VPWR _3597_ _4067_ _3133_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_89 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_1_120 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5373_ VPWR VGND _0683_ _0842_ _0841_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_8161_ VGND VPWR _3535_ _3064_ _3534_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_175 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7112_ VGND VPWR VPWR VGND _2561_ _2555_ _2563_ _1277_ _2562_ ZI_sky130_fd_sc_hd__o211a_2
X_8092_ VGND VPWR _3472_ _2640_ _3471_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4324_ VGND VPWR _3862_ _3861_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_112_489 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7043_ VGND VPWR VPWR VGND _2493_ _2485_ _2495_ _1277_ _2494_ ZI_sky130_fd_sc_hd__o211a_2
X_4255_ VGND VPWR VGND VPWR _3788_ _3789_ _3790_ _3791_ _3793_ _3792_ ZI_sky130_fd_sc_hd__o41ai_2
X_7945_ VGND VPWR _3339_ _4085_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_89_281 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7876_ VPWR VGND VPWR VGND _3219_ _3257_ _3276_ _3237_ _0801_ _3277_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_92_413 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6827_ VGND VPWR _2281_ _2280_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_65_627 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6758_ VPWR VGND _2139_ _2212_ _2175_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5709_ VPWR VGND VPWR VGND _1169_ _1173_ _1171_ _0708_ _1174_ ZI_sky130_fd_sc_hd__or4_2
X_6689_ VPWR VGND _2105_ _2143_ _2138_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_8428_ VGND VPWR VPWR VGND clk _0030_ reset_n new_block[115] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_579 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_103_445 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8359_ VGND VPWR VGND VPWR _3713_ _0444_ _3710_ _3711_ _3714_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_13_281 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_34_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5991_ VPWR VGND VGND VPWR _1436_ _1453_ _1349_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_91_57 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7730_ VPWR VGND _3144_ _1580_ _1565_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4942_ VPWR VGND VPWR VGND _0414_ _0413_ _0256_ _0286_ _0415_ ZI_sky130_fd_sc_hd__or4bb_2
X_7661_ VPWR VGND VPWR VGND _2796_ _4093_ _3080_ _2702_ _0238_ _3081_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_46_126 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_46_148 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6612_ sword_ctr_reg\[1\] _2066_ sword_ctr_reg\[0\] new_block[31] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
X_4873_ VGND VPWR VGND VPWR _3871_ _4021_ _3849_ _3983_ _0347_ ZI_sky130_fd_sc_hd__o22a_2
X_7592_ VPWR VGND VPWR VGND _2796_ _4093_ _3017_ _1909_ _0373_ _3018_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_40_72 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6543_ VGND VPWR _1999_ _1997_ _1998_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6474_ VPWR VGND VGND VPWR _1931_ _1861_ _1871_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_42_354 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_42_365 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_70_641 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5425_ VGND VPWR VGND VPWR _0894_ _0615_ _0670_ _0613_ ZI_sky130_fd_sc_hd__o21a_2
X_8213_ VGND VPWR VGND VPWR _3582_ _3581_ _3580_ _3579_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_2_473 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_112_253 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5356_ VPWR VGND _0591_ _0825_ _0639_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_8144_ VPWR VGND VGND VPWR _1563_ _3520_ _4089_ ZI_sky130_fd_sc_hd__nor2_2
X_5287_ VGND VPWR _0757_ _0635_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4307_ VPWR VGND VGND VPWR _3824_ _3831_ _3838_ _3844_ _3845_ ZI_sky130_fd_sc_hd__and4b_2
X_8075_ VPWR VGND _3457_ block[96] round_key[96] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7026_ _2228_ _2478_ _2126_ _2208_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_4238_ VGND VPWR VPWR VGND round[0] _3758_ _3779_ _3780_ ZI_sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_21_Right_21 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7928_ VGND VPWR _3323_ _3321_ _3322_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_92_210 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7859_ VPWR VGND _3261_ _2628_ _2552_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_108_526 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_52_118 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_30_Right_30 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_33_398 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_45_28 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_61_16 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_44_619 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_64_490 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_3_237 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_10_53 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_24_365 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5210_ VGND VPWR VGND VPWR _0680_ _0667_ _0662_ _0673_ _0679_ ZI_sky130_fd_sc_hd__a211o_2
X_6190_ VPWR VGND VGND VPWR _1651_ _1649_ _1650_ ZI_sky130_fd_sc_hd__nand2_2
X_5141_ VPWR VGND VPWR VGND _0610_ _0607_ _0602_ _0589_ _0597_ _0611_ ZI_sky130_fd_sc_hd__a221o_2
X_5072_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[107] sword_ctr_reg\[0\] _0542_
+ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_35_50 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5974_ VGND VPWR _1436_ _1435_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7713_ VGND VPWR VGND VPWR _3129_ _3128_ _3127_ _3126_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_59_273 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_19_137 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4925_ VGND VPWR VGND VPWR _4001_ _0398_ _0290_ _0395_ _0397_ ZI_sky130_fd_sc_hd__nand4b_2
X_4856_ VPWR VGND VGND VPWR _4181_ _3862_ _3955_ _3974_ _0330_ _0329_ ZI_sky130_fd_sc_hd__o221a_2
X_7644_ VPWR VGND _3065_ _3064_ _3054_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7575_ VGND VPWR _3002_ _2551_ _2639_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_181 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6526_ VPWR VGND VPWR VGND _1979_ _1981_ _1980_ _1978_ _1982_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_105_529 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4787_ VGND VPWR VGND VPWR _4003_ _4189_ _0183_ _0211_ _0262_ _0261_ ZI_sky130_fd_sc_hd__a2111o_2
X_6457_ VPWR VGND VPWR VGND _1592_ _1725_ _1602_ _1590_ _1914_ ZI_sky130_fd_sc_hd__or4_2
X_6388_ VPWR VGND VPWR VGND _1627_ _1845_ _1844_ _1598_ _1846_ ZI_sky130_fd_sc_hd__or4_2
X_5408_ VGND VPWR VGND VPWR _0877_ _0609_ _0605_ _0600_ _0598_ ZI_sky130_fd_sc_hd__and4_2
X_5339_ VPWR VGND _0809_ round_key[48] new_block[48] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8127_ VGND VPWR _3504_ _3009_ _3503_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8058_ VGND VPWR VGND VPWR _3441_ _0365_ _0811_ _4090_ _3442_ ZI_sky130_fd_sc_hd__a2bb2o_2
X_7009_ VPWR VGND VGND VPWR _2326_ _2461_ _2339_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_18_170 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_34_641 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_56_49 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4710_ VPWR VGND VGND VPWR _0186_ _3881_ _0185_ ZI_sky130_fd_sc_hd__nand2_2
X_5690_ VGND VPWR VGND VPWR _0757_ _0613_ _1154_ _0685_ _1155_ _0624_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_16_118 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4641_ VGND VPWR VPWR VGND _3898_ _3932_ _3857_ _4178_ ZI_sky130_fd_sc_hd__or3_2
X_7360_ VGND VPWR _2805_ _2802_ _2804_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_302 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_25_663 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4572_ VGND VPWR VPWR VGND _3891_ _3915_ _3831_ _4109_ ZI_sky130_fd_sc_hd__or3_2
X_6311_ VPWR VGND VPWR VGND _1281_ _0524_ _1770_ _0816_ _1769_ _1771_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_40_633 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7291_ VGND VPWR _2739_ _1146_ _2695_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6242_ VGND VPWR VPWR VGND _1700_ _1701_ _1594_ _1702_ ZI_sky130_fd_sc_hd__or3_2
X_6173_ VPWR VGND VPWR VGND _1631_ _1633_ _1634_ _1444_ _1462_ ZI_sky130_fd_sc_hd__or4b_2
X_5124_ VGND VPWR VPWR VGND _0574_ _0573_ _0572_ _4097_ _0575_ _0594_ ZI_sky130_fd_sc_hd__a41oi_2
X_5055_ VGND VPWR VGND VPWR _4104_ new_block[103] _0525_ _0521_ _0513_ _0018_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_27_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_122 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_1_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5957_ VGND VPWR _1419_ _1418_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4908_ VPWR VGND _0382_ round_key[92] new_block[92] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5888_ VPWR VGND VGND VPWR _1307_ _1350_ _1349_ ZI_sky130_fd_sc_hd__nor2_2
X_7627_ VGND VPWR VPWR VGND _3048_ _3046_ _3050_ _2855_ _3049_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_7_362 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_35_449 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4839_ VGND VPWR _0314_ _0310_ _0313_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7558_ VGND VPWR VGND VPWR _2894_ new_block[81] _2986_ _2983_ _1675_ _0060_ ZI_sky130_fd_sc_hd__o32a_2
X_6509_ VGND VPWR VGND VPWR _1940_ _1521_ _1390_ _1635_ _1965_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_15_195 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_30_121 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7489_ VPWR VGND VPWR VGND _2892_ _2786_ _2923_ _2880_ _0311_ _2924_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_97_165 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_42_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_109_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_66_585 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_53_246 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_108_153 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_108_197 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_6_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_21_176 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_83_69 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_16_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6860_ VPWR VGND _2314_ _2313_ _0818_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_88_165 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5811_ VGND VPWR _1274_ _1272_ _1273_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6791_ VPWR VGND _2182_ _2245_ _2070_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5742_ VGND VPWR VGND VPWR _1206_ _0678_ _0696_ _0664_ ZI_sky130_fd_sc_hd__o21a_2
X_8530_ VGND VPWR VPWR VGND clk _0132_ reset_n new_block[25] ZI_sky130_fd_sc_hd__dfrtp_2
X_5673_ VGND VPWR _1139_ _0799_ _1138_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8461_ VGND VPWR VPWR VGND clk _0063_ reset_n new_block[84] ZI_sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_6_Right_6 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_13_600 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7412_ VGND VPWR _2853_ _2851_ _2852_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4624_ VPWR VGND VGND VPWR _4159_ _4160_ _4161_ ZI_sky130_fd_sc_hd__or2b_2
X_8392_ VPWR VGND _3743_ _3191_ _1899_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7343_ VGND VPWR _2789_ _0904_ _2788_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4555_ VGND VPWR _4093_ _4092_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4486_ VGND VPWR VGND VPWR _4023_ _4021_ _4024_ _3990_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_110_340 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7274_ VPWR VGND VPWR VGND _2456_ _2101_ _2164_ _2131_ _2157_ _2722_ ZI_sky130_fd_sc_hd__a221o_2
X_6225_ VGND VPWR _1686_ _1682_ _1685_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6156_ VPWR VGND VPWR VGND _1471_ _1493_ _1523_ _1528_ _1617_ ZI_sky130_fd_sc_hd__a22o_2
X_5107_ VPWR VGND VGND VPWR _0576_ _0577_ _3880_ ZI_sky130_fd_sc_hd__nor2_2
X_6087_ VGND VPWR _1549_ _1548_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_79_143 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5038_ VGND VPWR VGND VPWR _3945_ _3949_ _3923_ _0509_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_48_541 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6989_ VGND VPWR VGND VPWR _2440_ _2128_ _2136_ _2297_ _2441_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_94_157 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_82_319 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_106_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_105_134 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_106_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_86_625 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_66_360 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_59_Right_59 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4340_ VGND VPWR _3878_ _3852_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4271_ VGND VPWR VGND VPWR _3797_ _3805_ _3806_ _3807_ _3809_ _3808_ ZI_sky130_fd_sc_hd__o41ai_2
X_6010_ VGND VPWR VPWR VGND _1318_ _1364_ _1312_ _1472_ ZI_sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_68_Right_68 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_27_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7961_ VGND VPWR VGND VPWR _3354_ _3353_ _3352_ _3348_ ZI_sky130_fd_sc_hd__o21a_2
X_7892_ VGND VPWR VGND VPWR _3291_ _3290_ _3289_ _2782_ ZI_sky130_fd_sc_hd__o21a_2
X_6912_ VPWR VGND VPWR VGND _2362_ _2364_ _2363_ _2360_ _2365_ ZI_sky130_fd_sc_hd__or4_2
X_6843_ VGND VPWR _2297_ _2138_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_43_83 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_99_Left_212 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6774_ VGND VPWR _2228_ _2227_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_77_Right_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_57_382 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_57_360 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5725_ VGND VPWR _1190_ _1187_ _1189_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8513_ VGND VPWR VPWR VGND clk _0115_ reset_n new_block[8] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5656_ VPWR VGND VPWR VGND _0889_ _1121_ _1120_ _0732_ _1122_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_94_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8444_ VGND VPWR VPWR VGND clk _0046_ reset_n new_block[67] ZI_sky130_fd_sc_hd__dfrtp_2
X_4607_ VGND VPWR VGND VPWR _4144_ _3959_ _4143_ _4142_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_32_249 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_102_126 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8375_ VGND VPWR VGND VPWR _3728_ _3727_ _3726_ _2944_ ZI_sky130_fd_sc_hd__o21a_2
X_5587_ VPWR VGND VPWR VGND _1040_ _1053_ _1045_ _1033_ _1054_ ZI_sky130_fd_sc_hd__or4_2
X_4538_ VPWR VGND _4076_ round_key[77] new_block[77] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7326_ VGND VPWR VPWR VGND _2767_ _2772_ _2334_ _2773_ ZI_sky130_fd_sc_hd__or3_2
X_7257_ VGND VPWR VGND VPWR _1911_ new_block[125] _2705_ _2701_ _2686_ _0040_ ZI_sky130_fd_sc_hd__o32a_2
X_4469_ VGND VPWR VPWR VGND _4004_ _4006_ _4001_ _4007_ ZI_sky130_fd_sc_hd__or3_2
X_6208_ VGND VPWR VGND VPWR _1669_ _1639_ _1456_ _1667_ _1668_ ZI_sky130_fd_sc_hd__a211o_2
XPHY_EDGE_ROW_86_Right_86 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_68_91 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7188_ VPWR VGND _2638_ _2637_ _2416_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6139_ VPWR VGND VPWR VGND _1332_ _1438_ _1379_ _1523_ _1600_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_68_625 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Right_95 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_83_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_55_308 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_63_374 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_90_193 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_63_396 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_23_249 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_59_625 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_59_658 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_74_628 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_27_522 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5510_ VGND VPWR VGND VPWR _0978_ _0639_ _0626_ _0698_ _0579_ ZI_sky130_fd_sc_hd__and4_2
XFILLER_0_109_281 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_27_599 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_89_57 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6490_ VGND VPWR _1947_ _1944_ _1946_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5441_ VPWR VGND _0910_ _0909_ _0798_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_89_68 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5372_ VGND VPWR _0841_ _0770_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8160_ VGND VPWR _3534_ _4064_ _0142_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7111_ VPWR VGND VGND VPWR _2562_ _2555_ _2561_ ZI_sky130_fd_sc_hd__nand2_2
X_8091_ VGND VPWR _3471_ _2421_ _2497_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4323_ VGND VPWR VPWR VGND _3852_ _3860_ _3794_ _3861_ ZI_sky130_fd_sc_hd__or3_2
X_7042_ VPWR VGND VGND VPWR _2494_ _2485_ _2493_ ZI_sky130_fd_sc_hd__nand2_2
X_4254_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[96] sword_ctr_reg\[0\] _3792_
+ ZI_sky130_fd_sc_hd__or3_2
X_7944_ VGND VPWR _3338_ _3335_ _3337_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_293 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7875_ VPWR VGND _3276_ block[109] round_key[109] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_49_135 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6826_ VPWR VGND _2070_ _2280_ _2133_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_65_639 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_18_533 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6757_ VGND VPWR VGND VPWR _2191_ _2128_ _2197_ _2198_ _2211_ _2210_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_92_447 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5708_ VPWR VGND VPWR VGND _1172_ _0628_ _0729_ _0602_ _0757_ _1173_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_70_81 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6688_ _2138_ _2142_ _2105_ _2141_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8427_ VGND VPWR VPWR VGND clk _0029_ reset_n new_block[114] ZI_sky130_fd_sc_hd__dfrtp_2
X_5639_ VGND VPWR VGND VPWR _0859_ _0616_ _0838_ _1102_ _1105_ _1104_ ZI_sky130_fd_sc_hd__a2111o_2
X_8358_ VPWR VGND VPWR VGND _3458_ _4093_ _3712_ _2702_ _1819_ _3713_ ZI_sky130_fd_sc_hd__a221o_2
X_7309_ VPWR VGND VPWR VGND _2752_ _2755_ _2753_ _2217_ _2756_ ZI_sky130_fd_sc_hd__or4_2
X_8289_ VGND VPWR VGND VPWR _3640_ new_block[20] _3650_ _3648_ _1884_ _0127_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_87_208 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_71_609 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_63_193 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_59_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5990_ VPWR VGND VGND VPWR _1368_ _1452_ _1307_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_99_580 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_78_219 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_24_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_59_455 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4941_ VPWR VGND VGND VPWR _3984_ _0414_ _3941_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_24_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_47_617 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7660_ VPWR VGND _3080_ block[90] round_key[90] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4872_ VPWR VGND VPWR VGND _4189_ _4168_ _3845_ _3926_ _0346_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_59_466 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_86_296 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6611_ VGND VPWR VGND VPWR _2065_ new_block[63] sword_ctr_reg\[1\] sword_ctr_reg\[0\]
+ ZI_sky130_fd_sc_hd__and3b_2
XFILLER_0_6_213 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7591_ VPWR VGND _3017_ block[116] round_key[116] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_39_190 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_6_246 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_6_257 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6542_ VGND VPWR _1998_ _1817_ _1833_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_82_491 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6473_ VPWR VGND VPWR VGND _1920_ _1929_ _1922_ _1916_ _1930_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_40_95 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5424_ VGND VPWR VGND VPWR _0893_ _0712_ _0666_ _0619_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_112_221 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8212_ VGND VPWR VGND VPWR _3580_ _3579_ _3581_ _3339_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_112_265 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8143_ VPWR VGND VPWR VGND _3519_ round_key[102] block[102] ZI_sky130_fd_sc_hd__or2_2
X_5355_ VPWR VGND VPWR VGND _0824_ _0822_ _0823_ ZI_sky130_fd_sc_hd__or2_2
XFILLER_0_57_3 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_10_274 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_10_296 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8074_ VGND VPWR VPWR VGND _3454_ _3452_ _3456_ _3448_ _3455_ ZI_sky130_fd_sc_hd__o211a_2
X_5286_ VGND VPWR VGND VPWR _0722_ _0754_ _0755_ _0756_ ZI_sky130_fd_sc_hd__a21o_2
X_4306_ VPWR VGND VGND VPWR _3844_ _3754_ _3843_ ZI_sky130_fd_sc_hd__nand2_2
X_7025_ _2166_ _2477_ _2297_ _2178_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_4237_ VPWR VGND VGND VPWR _3758_ _3779_ _0000_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_4_95 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7927_ VGND VPWR _3322_ _0231_ _0311_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7858_ VPWR VGND _3260_ _2639_ _2634_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_37_138 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6809_ VGND VPWR VGND VPWR _2263_ _2259_ _2107_ _2261_ _2262_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_92_222 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7789_ VGND VPWR VPWR VGND _3196_ _3195_ _3198_ _3118_ _3197_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_33_311 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_80_428 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Left_149 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_73_491 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_61_664 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_60_141 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_103_232 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Left_158 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_29_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_83_200 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_56_403 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_37_661 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_83_255 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_54_Left_167 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_24_322 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_52_631 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5140_ _0609_ _0610_ _0583_ _0592_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5071_ VGND VPWR VPWR VGND sword_ctr_reg\[0\] _0541_ new_block[43] ZI_sky130_fd_sc_hd__and2b_2
XPHY_EDGE_ROW_63_Left_176 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5973_ VGND VPWR VPWR VGND _1333_ _1392_ _3787_ _1435_ ZI_sky130_fd_sc_hd__or3_2
X_4924_ VPWR VGND VGND VPWR _0393_ _4181_ _3988_ _3955_ _0397_ _0396_ ZI_sky130_fd_sc_hd__o221a_2
X_7712_ VGND VPWR VGND VPWR _3127_ _3126_ _3128_ _3028_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_19_149 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4855_ VGND VPWR VGND VPWR _4131_ _3987_ _3984_ _0329_ ZI_sky130_fd_sc_hd__a21o_2
X_7643_ VGND VPWR _3064_ _0230_ _0435_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_72_Left_185 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_15_300 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7574_ VGND VPWR _3001_ _2491_ _3000_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4786_ VPWR VGND VGND VPWR _4025_ _0261_ _3887_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_74_277 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6525_ _1344_ _1981_ _1444_ _1379_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_55_491 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_42_141 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6456_ VPWR VGND VPWR VGND _1913_ _1454_ _1468_ ZI_sky130_fd_sc_hd__or2_2
X_6387_ VPWR VGND VPWR VGND _1424_ _1536_ _1341_ _1346_ _1845_ ZI_sky130_fd_sc_hd__a22o_2
X_5407_ VPWR VGND VPWR VGND _0864_ _0875_ _0869_ _0863_ _0876_ ZI_sky130_fd_sc_hd__or4_2
X_5338_ VGND VPWR _0808_ new_block[53] round_key[53] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8126_ VGND VPWR _3503_ _2693_ _3502_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_246 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_81_Left_194 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8057_ VGND VPWR _3441_ _2860_ _3440_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5269_ VPWR VGND _0557_ _0739_ _0608_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_7008_ VPWR VGND VPWR VGND _2434_ _2459_ _2446_ _2429_ _2460_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_76_80 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_80_214 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4640_ VPWR VGND VGND VPWR _3984_ _4114_ _4175_ _3982_ _4177_ _4176_ ZI_sky130_fd_sc_hd__o221a_2
X_6310_ VPWR VGND _1770_ new_block[114] round_key[114] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4571_ VGND VPWR VGND VPWR _4107_ _3894_ _3804_ _4030_ _4108_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_40_645 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7290_ VGND VPWR _2738_ _2310_ _2547_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6241_ VPWR VGND VPWR VGND _1499_ _1437_ _1331_ _1408_ _1701_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_97_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_110_533 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6172_ VPWR VGND VGND VPWR _1355_ _1531_ _1633_ _1381_ _1632_ ZI_sky130_fd_sc_hd__o22ai_2
X_5123_ VGND VPWR VGND VPWR _0593_ _4097_ _0526_ _0527_ _0528_ _0529_ ZI_sky130_fd_sc_hd__a41o_2
XFILLER_0_46_50 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5054_ VPWR VGND VPWR VGND _4101_ _0524_ _0523_ _0162_ _0522_ _0525_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_46_94 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5956_ _1318_ _1418_ _1352_ _1414_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5887_ VGND VPWR VPWR VGND _1347_ _1348_ _3796_ _1349_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_35_406 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4907_ VGND VPWR _0381_ _4073_ _0380_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7626_ VPWR VGND VGND VPWR _3049_ _3046_ _3048_ ZI_sky130_fd_sc_hd__nand2_2
X_4838_ VPWR VGND _0313_ _0312_ _4078_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_16_620 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_62_236 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7557_ VPWR VGND VPWR VGND _2892_ _2960_ _2985_ _2984_ _0152_ _2986_ ZI_sky130_fd_sc_hd__a221o_2
X_4769_ VGND VPWR _0245_ _0240_ _0244_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6508_ VPWR VGND VPWR VGND _1722_ _1776_ _1963_ _1494_ _1964_ ZI_sky130_fd_sc_hd__or4_2
X_7488_ VPWR VGND _2923_ block[11] round_key[11] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6439_ VPWR VGND _1897_ _1896_ _1895_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8109_ VGND VPWR VPWR VGND _3486_ _3485_ _3488_ _3448_ _3487_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_87_90 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_98_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_98_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_93_350 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_108_121 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_108_165 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_22_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_34_450 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_21_100 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_22_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_67_16 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_83_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_16_53 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_88_133 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_49_509 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5810_ VPWR VGND _1273_ _1126_ _0993_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_9_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6790_ VPWR VGND _2233_ _2244_ _2216_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_57_531 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_57_520 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5741_ VGND VPWR VGND VPWR _1205_ _0658_ _0635_ _0645_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_57_564 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8460_ VGND VPWR VPWR VGND clk _0062_ reset_n new_block[83] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_406 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_32_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5672_ VPWR VGND _1138_ round_key[43] new_block[43] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7411_ VGND VPWR _2852_ _0987_ _1133_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_85 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4623_ VGND VPWR VGND VPWR _4125_ _3971_ _3859_ _3992_ _4160_ ZI_sky130_fd_sc_hd__o22a_2
X_8391_ VPWR VGND _3742_ _3204_ _2003_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_72_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7342_ VPWR VGND _2788_ _0902_ _0807_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_13_612 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4554_ dec_ctrl_reg\[2\] _4092_ _3749_ _3766_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_40_453 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7273_ VGND VPWR VGND VPWR _2198_ _2163_ _2478_ _2209_ _2721_ _2720_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_12_177 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_40_497 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4485_ VGND VPWR _4023_ _4022_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6224_ VGND VPWR _1685_ _1683_ _1684_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6155_ VGND VPWR _1616_ _1493_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6086_ VGND VPWR VPWR VGND _1363_ _1398_ _1313_ _1548_ ZI_sky130_fd_sc_hd__or3_2
X_5106_ VGND VPWR VGND VPWR _0576_ _3828_ _0572_ _0573_ _0574_ _0575_ ZI_sky130_fd_sc_hd__a41o_2
X_5037_ VGND VPWR VGND VPWR _3981_ _3898_ _0503_ _0505_ _0508_ _0507_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_79_155 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_73_81 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6988_ VPWR VGND VPWR VGND _2186_ _2300_ _2190_ _2102_ _2440_ ZI_sky130_fd_sc_hd__a22o_2
X_5939_ VPWR VGND VGND VPWR _1401_ _1400_ _1369_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_75_350 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_63_501 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7609_ VGND VPWR _3033_ _1908_ _1961_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_113 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_106_625 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_86_637 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_85_103 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_39_553 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_39_575 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_54_567 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_112_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_111_105 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4270_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[98] sword_ctr_reg\[0\] _3808_
+ ZI_sky130_fd_sc_hd__or3_2
X_7960_ VGND VPWR VGND VPWR _3352_ _3348_ _3353_ _3339_ ZI_sky130_fd_sc_hd__a21oi_2
X_7891_ VGND VPWR VGND VPWR _3289_ _2782_ _3290_ _3028_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_89_475 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6911_ VPWR VGND VPWR VGND _2176_ _2167_ _2072_ _2106_ _2364_ ZI_sky130_fd_sc_hd__a22o_2
X_6842_ VPWR VGND _2112_ _2296_ _2212_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_43_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_43_73 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_9_436 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_91_106 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6773_ VPWR VGND VGND VPWR _2146_ _2227_ _2118_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_64_309 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5724_ VGND VPWR _1189_ _0995_ _1188_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_214 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_45_545 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8512_ VGND VPWR VPWR VGND clk _0114_ reset_n new_block[7] ZI_sky130_fd_sc_hd__dfrtp_2
X_5655_ VGND VPWR VGND VPWR _1121_ _0615_ _0612_ _0785_ _0975_ _0674_ ZI_sky130_fd_sc_hd__a32o_2
X_8443_ VGND VPWR VPWR VGND clk _0045_ reset_n new_block[66] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_5_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_87_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8374_ VGND VPWR VGND VPWR _3726_ _2944_ _3727_ _4085_ ZI_sky130_fd_sc_hd__a21oi_2
X_4606_ VPWR VGND VGND VPWR _4110_ _4143_ _3851_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_4_174 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_25_291 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_103_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7325_ VPWR VGND VPWR VGND _2769_ _2771_ _2770_ _2768_ _2772_ ZI_sky130_fd_sc_hd__or4_2
X_5586_ VPWR VGND VPWR VGND _0890_ _1052_ _1048_ _0759_ _1053_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_7_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4537_ VPWR VGND _4075_ round_key[80] new_block[80] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_102_149 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7256_ VPWR VGND VPWR VGND _4100_ _1959_ _2704_ _2703_ _2310_ _2705_ ZI_sky130_fd_sc_hd__a221o_2
X_4468_ _3903_ _4006_ _3795_ _4005_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6207_ VPWR VGND VPWR VGND _1476_ _1639_ _1421_ _1346_ _1522_ _1668_ ZI_sky130_fd_sc_hd__a221o_2
X_7187_ VPWR VGND _2637_ _0447_ _0363_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6138_ VGND VPWR VGND VPWR _1438_ _1340_ _1597_ _1598_ _1599_ _1402_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_110_193 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4399_ VGND VPWR VGND VPWR _3913_ _3911_ _3928_ _3931_ _3937_ _3936_ ZI_sky130_fd_sc_hd__a2111o_2
X_6069_ VGND VPWR _1531_ _1530_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_84_80 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_68_637 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_95_445 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_67_136 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_83_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_36_545 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_36_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_58_103 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_80_16 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_27_545 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_42_504 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5440_ VPWR VGND _0909_ _0908_ _0907_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_2_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_42_559 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_1_133 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_2_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5371_ VGND VPWR VPWR VGND _0838_ _0839_ _0646_ _0840_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_10_434 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7110_ VPWR VGND _2561_ _2560_ _2559_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4322_ VPWR VGND VPWR VGND _3814_ _3860_ _3787_ _3809_ ZI_sky130_fd_sc_hd__or3b_2
X_8090_ VGND VPWR VGND VPWR _3462_ new_block[1] _3470_ _3467_ _0140_ _0108_ ZI_sky130_fd_sc_hd__o32a_2
X_7041_ VGND VPWR _2493_ _2489_ _2492_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4253_ VGND VPWR VPWR VGND sword_ctr_reg\[0\] _3791_ new_block[32] ZI_sky130_fd_sc_hd__and2b_2
X_7943_ VGND VPWR _3337_ _0381_ _3336_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7874_ VGND VPWR VPWR VGND _3273_ _3272_ _3275_ _3265_ _3274_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_49_169 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6825_ VGND VPWR _2279_ _2278_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6756_ VGND VPWR VGND VPWR _2210_ _2178_ _2202_ _2206_ _2209_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_18_578 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5707_ VGND VPWR VGND VPWR _1172_ _0825_ _0684_ _0571_ _0729_ _0887_ ZI_sky130_fd_sc_hd__a32o_2
X_6687_ VGND VPWR _2141_ _2140_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8426_ VGND VPWR VPWR VGND clk _0028_ reset_n new_block[113] ZI_sky130_fd_sc_hd__dfrtp_2
X_5638_ VPWR VGND VPWR VGND _0628_ _0929_ _0602_ _1103_ _1104_ ZI_sky130_fd_sc_hd__a22o_2
X_8357_ VPWR VGND _3712_ block[27] round_key[27] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5569_ VGND VPWR VGND VPWR _0837_ _0724_ _0635_ _1036_ _0633_ ZI_sky130_fd_sc_hd__o2bb2a_2
X_7308_ VGND VPWR VGND VPWR _2755_ _2144_ _2136_ _2754_ _2108_ ZI_sky130_fd_sc_hd__a211o_2
X_8288_ VPWR VGND VPWR VGND _3575_ _3603_ _3649_ _3583_ _1945_ _3650_ ZI_sky130_fd_sc_hd__a221o_2
X_7239_ VGND VPWR _2688_ _2557_ _2687_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_180 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_63_161 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_91_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_99_592 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4940_ VGND VPWR VGND VPWR _0413_ _4189_ _3900_ _3845_ _4013_ _3795_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_24_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_86_253 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4871_ _3997_ _0345_ _3795_ _4134_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_24_97 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7590_ VGND VPWR _3016_ _3008_ _3015_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6610_ VPWR VGND VPWR VGND _2064_ new_block[126] _3828_ ZI_sky130_fd_sc_hd__or2_2
X_6541_ VPWR VGND _1997_ _1689_ _1578_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_55_640 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_27_375 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_6_269 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6472_ VGND VPWR VPWR VGND _1556_ _1928_ _1533_ _1929_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_40_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5423_ VGND VPWR VGND VPWR _0615_ _0690_ _0891_ _0741_ _0892_ ZI_sky130_fd_sc_hd__o22a_2
X_8211_ VGND VPWR _3580_ _0306_ _0517_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5354_ VPWR VGND VPWR VGND _0747_ _0771_ _0662_ _0658_ _0823_ ZI_sky130_fd_sc_hd__a22o_2
X_8142_ VPWR VGND VGND VPWR _3518_ round_key[102] block[102] ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_10_253 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_112_277 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4305_ VGND VPWR VGND VPWR _3797_ _3839_ _3840_ _3841_ _3842_ _3843_ ZI_sky130_fd_sc_hd__o41a_2
X_8073_ VPWR VGND VGND VPWR _3455_ _3452_ _3454_ ZI_sky130_fd_sc_hd__nand2_2
X_5285_ VPWR VGND VPWR VGND _0705_ _0639_ _0596_ _0544_ _0755_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_4_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7024_ VPWR VGND VGND VPWR _2476_ _2250_ _2475_ ZI_sky130_fd_sc_hd__nand2_2
X_4236_ VGND VPWR VGND VPWR _3768_ sword_ctr_reg\[1\] _3778_ _0006_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_4_85 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_69_209 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7926_ VGND VPWR _3321_ _4078_ _3073_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7857_ VGND VPWR _3259_ _2417_ _3038_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_81_81 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6808_ VPWR VGND VPWR VGND _2235_ _2260_ _2112_ _2255_ _2262_ ZI_sky130_fd_sc_hd__a22o_2
X_7788_ VPWR VGND VGND VPWR _3197_ _3195_ _3196_ ZI_sky130_fd_sc_hd__nand2_2
X_6739_ VPWR VGND VGND VPWR _2192_ _2193_ _2110_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_73_470 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_61_643 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8409_ VGND VPWR VPWR VGND clk _0011_ reset_n new_block[96] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_153 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_103_244 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_60_197 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_100_Left_213 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_88_529 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_29_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_36_161 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_3_217 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_107_561 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_51_142 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_101_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_86_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5070_ sword_ctr_reg\[1\] _0540_ sword_ctr_reg\[0\] new_block[11] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
X_5972_ VGND VPWR _1434_ _1433_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4923_ VGND VPWR VGND VPWR _3896_ _4115_ _4192_ _4131_ _0396_ ZI_sky130_fd_sc_hd__o22a_2
X_7711_ VPWR VGND _3127_ _0368_ _4067_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_87_551 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4854_ VPWR VGND VGND VPWR _4131_ _3993_ _3954_ _4114_ _0328_ _0327_ ZI_sky130_fd_sc_hd__o221a_2
X_7642_ VGND VPWR VGND VPWR _2997_ new_block[88] _3063_ _3061_ _2307_ _0067_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_15_312 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7573_ VPWR VGND _3000_ _2999_ _2317_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4785_ VPWR VGND VPWR VGND _4024_ _4055_ _4053_ _4004_ _0260_ ZI_sky130_fd_sc_hd__or4_2
X_6524_ VGND VPWR VGND VPWR _1980_ _1419_ _1501_ _1470_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_42_153 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_70_462 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6455_ VGND VPWR VGND VPWR _1912_ _1351_ _1355_ _1372_ _1539_ ZI_sky130_fd_sc_hd__a211o_2
X_6386_ VGND VPWR VGND VPWR _1527_ _1340_ _1514_ _1629_ _1844_ _1843_ ZI_sky130_fd_sc_hd__a2111o_2
X_5406_ VPWR VGND VPWR VGND _0871_ _0874_ _0872_ _0870_ _0875_ ZI_sky130_fd_sc_hd__or4_2
X_5337_ VPWR VGND _0807_ _0806_ _0805_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8125_ VGND VPWR _3502_ _2315_ _2633_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8056_ VGND VPWR _3440_ _3436_ _3439_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5268_ VGND VPWR VGND VPWR _0738_ _0656_ _0580_ _0666_ _0678_ _0704_ ZI_sky130_fd_sc_hd__a32o_2
X_7007_ VPWR VGND VPWR VGND _2451_ _2458_ _2453_ _2449_ _2459_ ZI_sky130_fd_sc_hd__or4_2
X_4219_ VGND VPWR VGND VPWR _3762_ _3764_ _3751_ dec_ctrl_reg\[0\] _3765_ ZI_sky130_fd_sc_hd__o22a_2
X_5199_ VGND VPWR _0669_ _0668_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7909_ VPWR VGND VGND VPWR _3306_ _3303_ _3305_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_65_256 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_80_226 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_0_209 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_96_392 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4570_ VGND VPWR VGND VPWR _4107_ _4105_ _3998_ _3930_ _4106_ ZI_sky130_fd_sc_hd__o211ai_2
XFILLER_0_52_451 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_52_462 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_108_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_24_164 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6240_ VPWR VGND _1613_ _1700_ _1426_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_40_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_110_501 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6171_ VPWR VGND VGND VPWR _1495_ _1632_ _1609_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_110_545 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5122_ VGND VPWR _0592_ _0591_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_110_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5053_ VGND VPWR _0524_ _0168_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_46_62 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_79_337 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5955_ VGND VPWR VGND VPWR _1412_ _1385_ _1417_ _1416_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_75_510 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5886_ VGND VPWR VGND VPWR _0538_ _1290_ _1291_ _1292_ _1293_ _1348_ ZI_sky130_fd_sc_hd__o41a_2
X_4906_ VGND VPWR _0380_ _0149_ _0234_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4837_ VGND VPWR _0312_ _0230_ _0311_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7625_ VGND VPWR _3048_ _2734_ _3047_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_120 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_16_632 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_62_248 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7556_ VPWR VGND _2985_ block[113] round_key[113] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4768_ VGND VPWR _0244_ _0242_ _0243_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6507_ VGND VPWR VPWR VGND _1963_ _1401_ _1384_ _1390_ _1737_ ZI_sky130_fd_sc_hd__o31ai_2
X_4699_ VGND VPWR VGND VPWR _0175_ _3949_ _0174_ _0173_ ZI_sky130_fd_sc_hd__o21a_2
X_7487_ VGND VPWR VPWR VGND _2920_ _2918_ _2922_ _2855_ _2921_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_70_270 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_31_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6438_ VGND VPWR _1896_ _1564_ _1831_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8108_ VPWR VGND VGND VPWR _3487_ _3485_ _3486_ ZI_sky130_fd_sc_hd__nand2_2
X_6369_ VGND VPWR _1828_ _1568_ _1570_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8039_ VGND VPWR _3424_ _1183_ _3423_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_613 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_97_123 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_98_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_34_462 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_108_177 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_22_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_22_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_83_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_88_112 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_8_106 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_9_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_29_245 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5740_ VGND VPWR VPWR VGND _1153_ _1203_ _1115_ _1204_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_57_554 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_32_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7410_ VGND VPWR _2851_ _2848_ _2850_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_546 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5671_ VPWR VGND _1137_ round_key[60] new_block[60] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8390_ VGND VPWR VGND VPWR _3461_ new_block[30] _3741_ _3739_ _2731_ _0137_ ZI_sky130_fd_sc_hd__o32a_2
X_4622_ _3939_ _4159_ _3869_ _4030_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_40_421 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4553_ VPWR VGND VGND VPWR _4081_ _4086_ _4091_ _4090_ _4087_ ZI_sky130_fd_sc_hd__o22ai_2
X_7341_ VGND VPWR VGND VPWR _4103_ new_block[127] _2787_ _2784_ _2775_ _0042_ ZI_sky130_fd_sc_hd__o32a_2
X_4484_ VPWR VGND VGND VPWR _4022_ _3881_ _3920_ ZI_sky130_fd_sc_hd__nand2_2
X_7272_ VPWR VGND _2345_ _2720_ _2265_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_6223_ VPWR VGND _1684_ round_key[1] new_block[1] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6154_ VPWR VGND VPWR VGND _1614_ _1527_ _1529_ _1337_ _1499_ _1615_ ZI_sky130_fd_sc_hd__a221o_2
X_5105_ VPWR VGND VGND VPWR sword_ctr_reg\[0\] sword_ctr_reg\[1\] new_block[104] _0575_
+ ZI_sky130_fd_sc_hd__nor3_2
X_6085_ VPWR VGND VGND VPWR _1547_ _1389_ _1381_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_32_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5036_ VPWR VGND VPWR VGND _0279_ _0506_ _0425_ _0174_ _0507_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_48_510 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6987_ VGND VPWR VGND VPWR _2439_ _2436_ _2118_ _2437_ _2438_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_73_93 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5938_ VPWR VGND VGND VPWR _1347_ _1400_ _3850_ ZI_sky130_fd_sc_hd__nor2_2
X_5869_ _1319_ _1331_ _1313_ _1330_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7608_ VGND VPWR VGND VPWR _2997_ new_block[85] _3032_ _3030_ _1943_ _0064_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_106_637 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7539_ VGND VPWR VGND VPWR _2894_ new_block[79] _2969_ _2967_ _1268_ _0058_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_43_281 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_101_331 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_94_660 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_26_215 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_93_181 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_112_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_94_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7890_ VGND VPWR _3289_ _3022_ _3288_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6910_ _2207_ _2363_ _2072_ _2162_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6841_ VPWR VGND _2084_ _2295_ _2294_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_9_404 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_76_137 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6772_ VPWR VGND VGND VPWR _2225_ _2226_ _2110_ ZI_sky130_fd_sc_hd__nor2_2
X_8511_ VGND VPWR VPWR VGND clk _0113_ reset_n new_block[6] ZI_sky130_fd_sc_hd__dfrtp_2
X_5723_ VPWR VGND _1188_ round_key[44] new_block[44] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_84_170 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5654_ VPWR VGND VPWR VGND _0601_ _0712_ _0690_ _0717_ _1120_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_45_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8442_ VGND VPWR VPWR VGND clk _0044_ reset_n new_block[65] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8373_ VPWR VGND _3726_ _3725_ _2938_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4605_ VPWR VGND VGND VPWR _4141_ _4142_ _3877_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_102_106 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_103_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7324_ VPWR VGND VPWR VGND _2177_ _2168_ _2072_ _2227_ _2771_ ZI_sky130_fd_sc_hd__a22o_2
X_5585_ VGND VPWR VPWR VGND _1050_ _1051_ _1049_ _1052_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_4_186 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4536_ VPWR VGND _4074_ _4073_ _4072_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7255_ VPWR VGND _2704_ block[125] round_key[125] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4467_ VPWR VGND VGND VPWR _3877_ _4005_ _3898_ ZI_sky130_fd_sc_hd__nor2_2
X_6206_ VPWR VGND VPWR VGND _1453_ _1531_ _1361_ _1438_ _1667_ ZI_sky130_fd_sc_hd__a22o_2
X_7186_ VGND VPWR _2636_ _2629_ _2635_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_110_161 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4398_ VGND VPWR _3935_ _3932_ _3936_ _3933_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
X_6137_ VPWR VGND VGND VPWR _1549_ _1598_ _1538_ ZI_sky130_fd_sc_hd__nor2_2
X_6068_ _1363_ _1530_ _1313_ _1414_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5019_ VGND VPWR VGND VPWR _4104_ new_block[102] _0490_ _0487_ _0475_ _0017_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_48_373 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_75_181 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_36_557 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_16_270 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_106_467 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_64_29 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_59_605 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_86_457 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_74_608 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_58_159 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_104_79 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_27_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_89_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_54_332 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_42_516 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_81_162 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_2_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_22_240 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5370_ VPWR VGND VPWR VGND _0746_ _0712_ _0546_ _0570_ _0839_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_22_273 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4321_ VGND VPWR _3859_ _3858_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7040_ VGND VPWR _2492_ _1006_ _2491_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4252_ sword_ctr_reg\[1\] _3790_ sword_ctr_reg\[0\] new_block[0] VPWR VGND VPWR VGND
+ ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_38_41 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7942_ VGND VPWR _3336_ _0312_ _0378_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_262 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7873_ VPWR VGND VGND VPWR _3274_ _3272_ _3273_ ZI_sky130_fd_sc_hd__nand2_2
X_6824_ VPWR VGND VGND VPWR _2192_ _2278_ _2095_ ZI_sky130_fd_sc_hd__nor2_2
X_6755_ _2203_ _2209_ _2207_ _2208_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5706_ VPWR VGND VPWR VGND _1170_ _0747_ _0702_ _0664_ _0661_ _1171_ ZI_sky130_fd_sc_hd__a221o_2
X_8425_ VGND VPWR VPWR VGND clk _0027_ reset_n new_block[112] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_505 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6686_ VPWR VGND _2133_ _2140_ _2139_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5637_ _0642_ _1103_ _0886_ _0643_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8356_ VPWR VGND VPWR VGND _3711_ _2920_ _3709_ ZI_sky130_fd_sc_hd__or2_2
X_5568_ VPWR VGND VPWR VGND _0771_ _0695_ _0747_ _0662_ _1035_ ZI_sky130_fd_sc_hd__a22o_2
X_8287_ VPWR VGND _3649_ block[52] round_key[52] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4519_ VPWR VGND VPWR VGND _4054_ _4056_ _4055_ _4053_ _4057_ ZI_sky130_fd_sc_hd__or4_2
X_7307_ VPWR VGND VPWR VGND _2190_ _2373_ _2345_ _2131_ _2754_ ZI_sky130_fd_sc_hd__a22o_2
X_5499_ VPWR VGND VPWR VGND _0607_ _0717_ _0664_ _0661_ _0967_ ZI_sky130_fd_sc_hd__a22o_2
X_7238_ VGND VPWR _2687_ _0250_ _0489_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7169_ VPWR VGND VPWR VGND _2373_ _2216_ _2327_ _2330_ _2619_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_95_221 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_49_660 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_48_192 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_76_490 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_91_471 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_91_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_24_65 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4870_ VPWR VGND VPWR VGND _4031_ _3913_ _3900_ _0185_ _0344_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_46_118 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6540_ VGND VPWR VPWR VGND _1996_ _1643_ _1973_ _1995_ _3755_ ZI_sky130_fd_sc_hd__o31a_2
XFILLER_0_55_652 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6471_ VPWR VGND VPWR VGND _1925_ _1927_ _1926_ _1923_ _1928_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_70_633 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_30_508 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5422_ VGND VPWR VGND VPWR _0891_ _0545_ _0596_ _0609_ _0698_ ZI_sky130_fd_sc_hd__and4_2
X_8210_ VGND VPWR _3579_ _3113_ _3578_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5353_ VPWR VGND VPWR VGND _0717_ _0740_ _0706_ _0689_ _0822_ ZI_sky130_fd_sc_hd__a22o_2
X_8141_ VGND VPWR VPWR VGND _3515_ _3510_ _3517_ _3448_ _3516_ ZI_sky130_fd_sc_hd__o211a_2
X_4304_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[102] sword_ctr_reg\[0\] _3842_
+ ZI_sky130_fd_sc_hd__or3_2
X_8072_ VGND VPWR _3454_ _2981_ _3453_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_84 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5284_ VPWR VGND VGND VPWR _0543_ _0754_ _3776_ ZI_sky130_fd_sc_hd__nor2_2
X_7023_ VGND VPWR VGND VPWR _2196_ _2372_ _2475_ _2395_ ZI_sky130_fd_sc_hd__a21oi_2
X_4235_ VGND VPWR VGND VPWR _3771_ _3770_ _3778_ _3777_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_4_53 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_65_83 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7925_ VPWR VGND _3320_ _3054_ _0302_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7856_ VGND VPWR VGND VPWR _3240_ new_block[43] _3258_ _3255_ _1054_ _0086_ ZI_sky130_fd_sc_hd__o32a_2
X_6807_ VPWR VGND _2167_ _2261_ _2260_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_4999_ VGND VPWR VGND VPWR _4016_ _3918_ _0471_ _3982_ ZI_sky130_fd_sc_hd__a21oi_2
X_7787_ VGND VPWR _3196_ _1895_ _1955_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_365 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6738_ VGND VPWR VGND VPWR _2083_ _2078_ _2192_ _3880_ ZI_sky130_fd_sc_hd__a21oi_2
X_6669_ VGND VPWR _2123_ _2122_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8408_ VGND VPWR VPWR VGND clk _0010_ reset_n round[3] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_292 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_103_267 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8339_ VPWR VGND VGND VPWR _3521_ _3695_ _0162_ _3693_ _3694_ _3696_ ZI_sky130_fd_sc_hd__a311o_2
XFILLER_0_24_302 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_52_611 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_51_121 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_107_573 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_51_154 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_20_585 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_35_31 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5971_ _1362_ _1433_ _1312_ _1330_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_4922_ VPWR VGND VGND VPWR _0393_ _4131_ _3984_ _3933_ _0395_ _0394_ ZI_sky130_fd_sc_hd__o221a_2
X_7710_ VGND VPWR _3126_ _3124_ _3125_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7641_ VPWR VGND VPWR VGND _2995_ _3062_ _2857_ _2984_ _4063_ _3063_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_28_641 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4853_ VGND VPWR VGND VPWR _3998_ _4115_ _3999_ _4021_ _0327_ ZI_sky130_fd_sc_hd__o22a_2
XFILLER_0_47_449 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_51_52 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_27_162 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7572_ VGND VPWR _2999_ _2412_ _2625_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_611 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4784_ VPWR VGND VPWR VGND _0255_ _0258_ _0257_ _0253_ _0259_ ZI_sky130_fd_sc_hd__or4_2
X_6523_ VPWR VGND VPWR VGND _1339_ _1456_ _1360_ _1470_ _1979_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_42_121 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6454_ VGND VPWR VGND VPWR _1911_ new_block[116] _1910_ _1906_ _1884_ _0031_ ZI_sky130_fd_sc_hd__o32a_2
X_5405_ VPWR VGND VPWR VGND _0873_ _0589_ _0696_ _0746_ _0645_ _0874_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_42_165 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6385_ VGND VPWR VGND VPWR _1843_ _1530_ _1381_ _1437_ _1489_ _1344_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_100_204 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5336_ VPWR VGND _0806_ round_key[56] new_block[56] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8124_ VGND VPWR VGND VPWR _3462_ new_block[4] _3501_ _3499_ _0362_ _0111_ ZI_sky130_fd_sc_hd__o32a_2
X_8055_ VGND VPWR _3439_ _3437_ _3438_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5267_ VGND VPWR VGND VPWR _0737_ _0571_ _0710_ _0671_ ZI_sky130_fd_sc_hd__o21a_2
X_4218_ VGND VPWR _3764_ _3763_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7006_ VGND VPWR VGND VPWR _2246_ _2336_ _2454_ _2455_ _2458_ _2457_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_76_93 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5198_ VPWR VGND _0586_ _0668_ _0568_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_92_81 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7908_ VGND VPWR _3305_ _3085_ _3304_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7839_ VGND VPWR _3243_ _0818_ _2552_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_235 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_34_611 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_108_348 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_65_268 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_88_305 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_72_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_69_541 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_29_405 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_29_449 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_84_533 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_44_408 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_4_505 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_52_430 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_112_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_97_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_110_513 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6170_ VGND VPWR VPWR VGND _1629_ _1630_ _1372_ _1631_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_110_557 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5121_ VPWR VGND VGND VPWR _3879_ _0537_ _0590_ _0591_ ZI_sky130_fd_sc_hd__nor3_2
XFILLER_0_46_41 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5052_ VPWR VGND _0523_ new_block[103] round_key[103] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_46_74 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5954_ VGND VPWR _1416_ _1415_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5885_ VGND VPWR VGND VPWR _0538_ _1283_ _1284_ _1285_ _1347_ _1286_ ZI_sky130_fd_sc_hd__o41ai_2
X_4905_ VPWR VGND _0379_ _0378_ _0375_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_87_393 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4836_ VPWR VGND _0311_ round_key[75] new_block[75] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7624_ VPWR VGND _3047_ _2557_ _0363_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7555_ VGND VPWR _2984_ _2702_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_15_132 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6506_ VGND VPWR VGND VPWR _1911_ new_block[117] _1962_ _1958_ _1943_ _0032_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_43_452 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4767_ VPWR VGND _0243_ _0147_ _0143_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_15_176 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4698_ VGND VPWR VGND VPWR _3913_ _3900_ _3853_ _3871_ _0174_ ZI_sky130_fd_sc_hd__a2bb2o_2
X_7486_ VPWR VGND VGND VPWR _2921_ _2918_ _2920_ ZI_sky130_fd_sc_hd__nand2_2
X_6437_ VPWR VGND _1895_ round_key[4] new_block[4] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6368_ VGND VPWR _1827_ _1823_ _1826_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8107_ VPWR VGND _3486_ _3230_ _2484_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5319_ VGND VPWR VGND VPWR _0787_ _0747_ _0788_ _0789_ ZI_sky130_fd_sc_hd__a21o_2
X_6299_ VPWR VGND _1759_ round_key[17] new_block[17] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8038_ VGND VPWR _3423_ _1128_ _2875_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_157 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_38_202 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_66_533 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_22_625 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_21_146 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_83_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_107_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5670_ VGND VPWR _1136_ _0901_ _1135_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_257 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_32_65 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_32_98 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4621_ VGND VPWR VGND VPWR _3987_ _3896_ _4158_ _3969_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_72_558 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4552_ VGND VPWR _4090_ _4089_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7340_ VPWR VGND VPWR VGND _4100_ _2786_ _2785_ _2703_ _2311_ _2787_ ZI_sky130_fd_sc_hd__a221o_2
X_4483_ VGND VPWR _4021_ _4020_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7271_ VGND VPWR VGND VPWR _2283_ _2219_ _2132_ _2282_ _2719_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_40_477 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6222_ VGND VPWR _1683_ new_block[7] round_key[7] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_574 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6153_ VPWR VGND _1613_ _1614_ _1409_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_57_62 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6084_ VPWR VGND VGND VPWR _1399_ _1546_ _1436_ ZI_sky130_fd_sc_hd__nor2_2
X_5104_ VGND VPWR VGND VPWR sword_ctr_reg\[1\] sword_ctr_reg\[0\] new_block[72] _0574_
+ ZI_sky130_fd_sc_hd__nand3b_2
X_5035_ VGND VPWR VGND VPWR _3961_ _3999_ _0506_ _3974_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_25_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_79_124 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_95_606 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_69_Left_182 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_95_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6986_ VPWR VGND VPWR VGND _2228_ _2300_ _2170_ _2177_ _2438_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_67_308 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5937_ VGND VPWR VPWR VGND _1319_ _1398_ _1353_ _1399_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_48_522 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_48_533 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7607_ VPWR VGND VPWR VGND _2995_ _3031_ _2857_ _2984_ _4072_ _3032_ ZI_sky130_fd_sc_hd__a221o_2
X_5868_ VPWR VGND VGND VPWR _3775_ _1330_ _1329_ _1324_ ZI_sky130_fd_sc_hd__nor3b_2
XFILLER_0_63_536 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_105_104 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4819_ VGND VPWR VPWR VGND _0274_ _0293_ _0264_ _0294_ ZI_sky130_fd_sc_hd__or3_2
X_5799_ VGND VPWR VGND VPWR _1262_ _0771_ _0765_ _0671_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_16_485 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7538_ VPWR VGND VPWR VGND _2892_ _2960_ _2968_ _2880_ _0230_ _2969_ ZI_sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_78_Left_191 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7469_ VGND VPWR _2905_ _2903_ _2904_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_591 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_19_Right_19 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_39_511 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_85_116 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_26_227 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_39_599 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_81_322 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_66_385 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_26_249 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_93_193 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_28_Right_28 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_27_76 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_27_98 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_37_Right_37 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_89_444 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_89_499 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6840_ _2138_ _2294_ _2252_ _2175_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_77_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_76_105 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6771_ VGND VPWR VGND VPWR _2182_ _2099_ _2225_ _2100_ ZI_sky130_fd_sc_hd__nand3_2
XFILLER_0_69_190 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5722_ VGND VPWR _1187_ _1185_ _1186_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8510_ VGND VPWR VPWR VGND clk _0112_ reset_n new_block[5] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_84_182 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_5_611 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5653_ VGND VPWR VPWR VGND _1117_ _1118_ _1116_ _1119_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_60_506 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8441_ VGND VPWR VPWR VGND clk _0043_ reset_n new_block[64] ZI_sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_46_Right_46 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8372_ VGND VPWR _3725_ _2927_ _3724_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_528 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4604_ VGND VPWR _4141_ _4140_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5584_ _0580_ _1051_ _0688_ _0785_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_13_444 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4535_ VPWR VGND _4073_ round_key[86] new_block[86] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7323_ VGND VPWR VGND VPWR _2770_ _2285_ _2158_ _2123_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_111_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7254_ VGND VPWR _2703_ _2702_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4466_ VPWR VGND VPWR VGND _3913_ _4003_ _4002_ _3950_ _4004_ ZI_sky130_fd_sc_hd__a22o_2
X_6205_ VPWR VGND VPWR VGND _1500_ _1665_ _1664_ _1417_ _1666_ ZI_sky130_fd_sc_hd__or4_2
X_7185_ VGND VPWR _2635_ _2631_ _2634_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_110_173 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4397_ VPWR VGND VGND VPWR _3935_ _3903_ _3934_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_0_393 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6136_ VPWR VGND VGND VPWR _1460_ _1597_ _1416_ ZI_sky130_fd_sc_hd__nor2_2
X_6067_ VGND VPWR _1529_ _1528_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_55_Right_55 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5018_ VPWR VGND VPWR VGND _4101_ _0169_ _0489_ _0162_ _0488_ _0490_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_67_105 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6969_ VPWR VGND VPWR VGND _4100_ _1909_ _2421_ _1959_ _2420_ _2422_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_82_108 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_36_569 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_91_642 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_75_193 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_63_388 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_16_293 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Right_73 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_80_29 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_67_650 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_27_514 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_82_Right_82 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_42_528 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_89_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_81_196 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_112_449 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4320_ VGND VPWR VPWR VGND _3857_ _3852_ _3851_ _3858_ ZI_sky130_fd_sc_hd__or3_2
X_4251_ VGND VPWR VGND VPWR _3789_ sword_ctr_reg\[0\] new_block[64] sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__and3b_2
XPHY_EDGE_ROW_91_Right_91 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_38_64 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7941_ VGND VPWR _3335_ _3333_ _3334_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7872_ VPWR VGND _3273_ _2692_ _2690_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_54_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6823_ VPWR VGND VPWR VGND _2263_ _2276_ _2270_ _2258_ _2277_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_65_609 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6754_ VGND VPWR _2208_ _2195_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5705_ VPWR VGND VPWR VGND _0651_ _0690_ _0545_ _0678_ _1170_ ZI_sky130_fd_sc_hd__a22o_2
X_6685_ VGND VPWR VGND VPWR _2139_ _2064_ _2063_ _2098_ _3753_ ZI_sky130_fd_sc_hd__and4_2
X_8424_ VGND VPWR VPWR VGND clk _0026_ reset_n new_block[111] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_92_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5636_ VGND VPWR VGND VPWR _1102_ _0616_ _0580_ _0669_ _0602_ _0674_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_41_561 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8355_ VPWR VGND VGND VPWR _3710_ _2920_ _3709_ ZI_sky130_fd_sc_hd__nand2_2
X_5567_ VGND VPWR VGND VPWR _1034_ _0975_ _0662_ _0706_ ZI_sky130_fd_sc_hd__o21a_2
X_8286_ VGND VPWR VGND VPWR _3648_ _3647_ _3646_ _3645_ ZI_sky130_fd_sc_hd__o21a_2
X_4518_ VGND VPWR VGND VPWR _4016_ _3983_ _4056_ _3992_ ZI_sky130_fd_sc_hd__a21oi_2
X_7306_ VGND VPWR VGND VPWR _2174_ _2327_ _2275_ _2753_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_79_93 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5498_ VPWR VGND VPWR VGND _0710_ _0648_ _0747_ _0589_ _0966_ ZI_sky130_fd_sc_hd__a22o_2
X_4449_ VGND VPWR _3987_ _3916_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7237_ VGND VPWR VPWR VGND _2663_ _2685_ _2657_ _2686_ ZI_sky130_fd_sc_hd__or3_2
X_7168_ VPWR VGND VPWR VGND _2618_ _2273_ ZI_sky130_fd_sc_hd__inv_2
X_7099_ VGND VPWR _2550_ _0818_ _2411_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6119_ VGND VPWR _1581_ _1577_ _1580_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_83_417 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_63_130 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_106_221 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_91_483 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_99_561 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_91_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_47_609 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_24_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_70_612 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6470_ VGND VPWR VGND VPWR _1927_ _1421_ _1353_ _1419_ _1471_ _1338_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_70_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5421_ VGND VPWR VPWR VGND _0885_ _0889_ _0884_ _0890_ ZI_sky130_fd_sc_hd__or3_2
X_5352_ VPWR VGND VPWR VGND _0820_ _0639_ _0761_ _0689_ _0787_ _0821_ ZI_sky130_fd_sc_hd__a221o_2
X_8140_ VPWR VGND VGND VPWR _3516_ _3510_ _3515_ ZI_sky130_fd_sc_hd__nand2_2
X_8071_ VGND VPWR _3453_ _0489_ _2011_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4303_ VGND VPWR VGND VPWR _3841_ sword_ctr_reg\[0\] new_block[70] sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__and3b_2
XFILLER_0_49_96 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7022_ VPWR VGND VPWR VGND _2474_ _2472_ _2473_ ZI_sky130_fd_sc_hd__or2_2
X_5283_ VPWR VGND VPWR VGND _0752_ _0753_ _0744_ _0750_ ZI_sky130_fd_sc_hd__or3b_2
X_4234_ VGND VPWR _3777_ _3776_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7924_ VGND VPWR VGND VPWR _3240_ new_block[50] _3319_ _3317_ _1750_ _0093_ ZI_sky130_fd_sc_hd__o32a_2
X_7855_ VPWR VGND VPWR VGND _3219_ _3257_ _3256_ _3237_ _1138_ _3258_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_77_233 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_46_620 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6806_ VGND VPWR _2260_ _2239_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_18_322 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7786_ VGND VPWR _3195_ _3192_ _3194_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4998_ VPWR VGND VPWR VGND _0469_ _0470_ _0339_ _0420_ ZI_sky130_fd_sc_hd__or3b_2
XFILLER_0_18_377 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6737_ VGND VPWR VGND VPWR _2191_ _2127_ _2073_ _2178_ _2190_ _2187_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_61_612 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_45_185 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6668_ VPWR VGND _2113_ _2122_ _2121_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_60_111 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_33_358 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8407_ VGND VPWR VPWR VGND clk _0009_ reset_n round[2] ZI_sky130_fd_sc_hd__dfrtp_2
X_6599_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[125] sword_ctr_reg\[0\] _2053_
+ ZI_sky130_fd_sc_hd__or3_2
X_5619_ VGND VPWR VGND VPWR _1084_ _0674_ _0689_ _0888_ _1085_ ZI_sky130_fd_sc_hd__a31o_2
X_8338_ VPWR VGND VGND VPWR _1679_ _3695_ _4089_ ZI_sky130_fd_sc_hd__nor2_2
X_8269_ VPWR VGND _3632_ _1071_ _0992_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_14_Left_127 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_29_609 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_36_141 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_36_185 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_52_623 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_52_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_101_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_107_541 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_107_585 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_136 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_51_188 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_108_Right_108 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5970_ VPWR VGND _1381_ _1432_ _1396_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_32_Left_145 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4921_ VGND VPWR VGND VPWR _4115_ _3976_ _3969_ _3885_ _3838_ _0394_ ZI_sky130_fd_sc_hd__o32a_2
X_4852_ VPWR VGND VGND VPWR _3962_ _4023_ _3999_ _4116_ _0326_ _0325_ ZI_sky130_fd_sc_hd__o221a_2
X_7640_ VPWR VGND _3062_ block[88] round_key[88] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_28_653 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_28_664 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7571_ VGND VPWR _2998_ _2416_ _2559_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4783_ VGND VPWR VGND VPWR _4105_ _3965_ _0258_ _4046_ ZI_sky130_fd_sc_hd__a21oi_2
X_6522_ VPWR VGND VPWR VGND _1613_ _1493_ _1394_ _1499_ _1978_ ZI_sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_41_Left_154 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_43_667 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6453_ VGND VPWR _1911_ _4103_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_30_328 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5404_ VGND VPWR VGND VPWR _0873_ _0596_ _0592_ _0609_ _0583_ ZI_sky130_fd_sc_hd__and4_2
X_6384_ VGND VPWR VGND VPWR _1009_ new_block[115] _1842_ _1839_ _1815_ _0030_ ZI_sky130_fd_sc_hd__o32a_2
X_8123_ VPWR VGND VPWR VGND _3459_ _3490_ _3500_ _3468_ _1895_ _3501_ ZI_sky130_fd_sc_hd__a221o_2
X_5335_ VGND VPWR _0805_ new_block[61] round_key[61] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8054_ VGND VPWR _3438_ _0913_ _1188_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5266_ _0705_ _0736_ _0583_ _0609_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_55_3 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4217_ VPWR VGND VPWR VGND _3763_ sword_ctr_reg\[1\] ZI_sky130_fd_sc_hd__inv_2
X_7005_ VPWR VGND _2163_ _2457_ _2456_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5197_ VPWR VGND VPWR VGND _0667_ _0664_ _0666_ ZI_sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_50_Left_163 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7907_ VGND VPWR _3304_ _0307_ _0386_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7838_ VGND VPWR _3242_ _3010_ _3241_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_19_653 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7769_ VGND VPWR VGND VPWR _3153_ new_block[35] _3179_ _3177_ _0294_ _0078_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_34_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_104_533 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_69_553 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_84_556 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_56_225 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_112_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_24_155 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_97_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_110_525 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_110_569 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5120_ VGND VPWR VGND VPWR _3788_ _0539_ _0540_ _0541_ _0542_ _0590_ ZI_sky130_fd_sc_hd__o41a_2
X_5051_ VPWR VGND _0522_ block[71] round_key[71] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_94_309 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5953_ VPWR VGND VPWR VGND _1414_ _1415_ _1312_ _1362_ ZI_sky130_fd_sc_hd__or3b_2
XFILLER_0_87_350 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5884_ VGND VPWR _1346_ _1345_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4904_ VGND VPWR _0378_ _0155_ _0377_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_450 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7623_ VGND VPWR _3046_ _3044_ _3045_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4835_ VPWR VGND _0310_ _0309_ _0307_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7554_ VGND VPWR VGND VPWR _2983_ _2982_ _2981_ _2980_ ZI_sky130_fd_sc_hd__o21a_2
X_4766_ VPWR VGND _0242_ _0241_ _4067_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_16_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6505_ VPWR VGND VPWR VGND _1281_ _1909_ _1961_ _1959_ _1960_ _1962_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_31_604 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4697_ VPWR VGND VGND VPWR _4125_ _0173_ _3933_ ZI_sky130_fd_sc_hd__nor2_2
X_7485_ VPWR VGND _2920_ _2919_ _1691_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6436_ VPWR VGND _1894_ _1752_ _1683_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_30_169 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6367_ VGND VPWR _1826_ _1824_ _1825_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8106_ VGND VPWR _3485_ _3483_ _3484_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5318_ VGND VPWR VGND VPWR _0788_ _0569_ _0591_ _0605_ _0598_ ZI_sky130_fd_sc_hd__and4_2
X_6298_ VGND VPWR _1758_ _1754_ _1757_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5249_ VGND VPWR VGND VPWR _0712_ _0710_ _0714_ _0715_ _0719_ _0718_ ZI_sky130_fd_sc_hd__a2111o_2
X_8037_ VGND VPWR VGND VPWR new_block[60] _3153_ _2624_ _3422_ _0103_ ZI_sky130_fd_sc_hd__o22a_2
XFILLER_0_97_169 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_66_512 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_38_214 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_66_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_22_637 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_21_158 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_107_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_29_225 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_29_269 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_57_578 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_32_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4620_ VGND VPWR VPWR VGND _4147_ _4156_ _4137_ _4157_ ZI_sky130_fd_sc_hd__or3_2
X_4551_ VGND VPWR _4089_ _4088_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4482_ VGND VPWR VPWR VGND _3852_ _3876_ _3794_ _4020_ ZI_sky130_fd_sc_hd__or3_2
X_7270_ VGND VPWR VPWR VGND _2715_ _2717_ _2357_ _2718_ ZI_sky130_fd_sc_hd__or3_2
X_6221_ VGND VPWR _1682_ _1574_ _1681_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6152_ VPWR VGND VGND VPWR _1307_ _1613_ _1389_ ZI_sky130_fd_sc_hd__nor2_2
X_5103_ VGND VPWR VGND VPWR sword_ctr_reg\[0\] new_block[40] sword_ctr_reg\[1\] _0573_
+ ZI_sky130_fd_sc_hd__nand3b_2
X_6083_ VGND VPWR VGND VPWR _1531_ _1395_ _1542_ _1543_ _1545_ _1544_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_57_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_57_74 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5034_ VGND VPWR VGND VPWR _0504_ _3967_ _3869_ _3925_ _0505_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_18_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6985_ VGND VPWR VGND VPWR _2437_ _2126_ _2072_ _2256_ _2302_ _2186_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_95_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5936_ VPWR VGND VPWR VGND _1324_ _1398_ _3850_ _1329_ ZI_sky130_fd_sc_hd__or3b_2
XFILLER_0_48_578 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_7_141 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7606_ VPWR VGND _3031_ block[117] round_key[117] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5867_ VGND VPWR VGND VPWR _3797_ _1325_ _1326_ _1327_ _1329_ _1328_ ZI_sky130_fd_sc_hd__o41ai_2
X_4818_ VPWR VGND VPWR VGND _0281_ _0292_ _0293_ _4113_ _0194_ ZI_sky130_fd_sc_hd__or4b_2
XFILLER_0_90_345 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5798_ VPWR VGND VPWR VGND _0958_ _0961_ _0960_ _0779_ _1261_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_63_548 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7537_ VPWR VGND _2968_ block[15] round_key[15] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4749_ VGND VPWR VGND VPWR _4031_ _4042_ _3941_ _3854_ _0225_ ZI_sky130_fd_sc_hd__a2bb2o_2
X_7468_ VPWR VGND _2904_ _1690_ _1579_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6419_ VPWR VGND _1340_ _1877_ _1604_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_7399_ VGND VPWR _2841_ _2834_ _2840_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_489 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_39_501 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_85_128 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_26_239 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_109_488 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_78_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_104_160 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_6_Left_119 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_27_88 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_77_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_43_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6770_ VPWR VGND _2222_ _2224_ _2223_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_76_117 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5721_ VPWR VGND _1186_ _0805_ _0808_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5652_ VGND VPWR VGND VPWR _1118_ _0888_ _0695_ _0664_ ZI_sky130_fd_sc_hd__o21a_2
X_8440_ VGND VPWR VPWR VGND clk _0042_ reset_n new_block[127] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_111 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8371_ VGND VPWR _3724_ _1886_ _3723_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_389 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4603_ VGND VPWR VPWR VGND _3838_ _3885_ _3831_ _4140_ ZI_sky130_fd_sc_hd__or3_2
X_5583_ VPWR VGND VPWR VGND _0664_ _0841_ _0627_ _0710_ _1050_ ZI_sky130_fd_sc_hd__a22o_2
X_4534_ VPWR VGND _4072_ round_key[85] new_block[85] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_53_581 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_103_609 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7322_ VPWR VGND VPWR VGND _2072_ _2279_ _2148_ _2213_ _2769_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_111_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4465_ VPWR VGND VGND VPWR _3910_ _4003_ _3932_ ZI_sky130_fd_sc_hd__nor2_2
X_7253_ VGND VPWR _2702_ _0168_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6204_ VGND VPWR VGND VPWR _1410_ _1534_ _1359_ _1616_ _1665_ ZI_sky130_fd_sc_hd__a31o_2
X_7184_ VGND VPWR _2634_ _2632_ _2633_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4396_ VPWR VGND VGND VPWR _3932_ _3934_ _3803_ ZI_sky130_fd_sc_hd__nor2_2
X_6135_ VGND VPWR VPWR VGND _1591_ _1595_ _1540_ _1596_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_110_185 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6066_ _1363_ _1528_ _1353_ _1330_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5017_ VPWR VGND _0489_ new_block[102] round_key[102] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6968_ VPWR VGND _2421_ new_block[121] round_key[121] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5919_ VGND VPWR _1381_ _1380_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6899_ VPWR VGND _2215_ _2352_ _2267_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_75_150 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_8_472 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_91_654 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_90_153 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_101_163 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_98_242 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_98_253 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_98_264 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_86_404 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_104_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_67_662 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_39_386 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_89_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_54_378 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_1_103 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_2_637 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_22_220 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_50_551 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4250_ VPWR VGND VGND VPWR sword_ctr_reg\[1\] _3788_ sword_ctr_reg\[0\] ZI_sky130_fd_sc_hd__nor2_2
X_7940_ VPWR VGND _3334_ _0386_ _0382_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7871_ VGND VPWR _3272_ _3270_ _3271_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_75 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_89_275 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6822_ VPWR VGND VPWR VGND _2272_ _2275_ _2274_ _2271_ _2276_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_9_203 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6753_ VPWR VGND VGND VPWR _2207_ _2118_ _2188_ ZI_sky130_fd_sc_hd__nand2_2
X_5704_ VPWR VGND VPWR VGND _1168_ _0748_ _0975_ _0675_ _0661_ _1169_ ZI_sky130_fd_sc_hd__a221o_2
X_6684_ VPWR VGND VGND VPWR _3775_ _2138_ _2094_ _2089_ ZI_sky130_fd_sc_hd__nor3b_2
XFILLER_0_72_131 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_70_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8423_ VGND VPWR VPWR VGND clk _0025_ reset_n new_block[110] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_72_153 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5635_ VGND VPWR VPWR VGND _0964_ _1100_ _0883_ _1101_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_60_304 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_85_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5566_ VPWR VGND VPWR VGND _1023_ _1032_ _1028_ _1017_ _1033_ ZI_sky130_fd_sc_hd__or4_2
X_8354_ VGND VPWR _3709_ _1835_ _3708_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8285_ VGND VPWR VGND VPWR _3646_ _3645_ _3647_ _4085_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_41_573 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7305_ VPWR VGND _2150_ _2752_ _2336_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5497_ VPWR VGND VPWR VGND _0964_ _0923_ _0963_ _0695_ _0748_ _0965_ ZI_sky130_fd_sc_hd__a221o_2
X_4517_ VGND VPWR VGND VPWR _3921_ _3918_ _4055_ _3872_ ZI_sky130_fd_sc_hd__a21oi_2
X_4448_ VPWR VGND VGND VPWR _3982_ _3986_ _3974_ ZI_sky130_fd_sc_hd__nor2_2
X_7236_ VPWR VGND VPWR VGND _2678_ _2684_ _2679_ _2670_ _2685_ ZI_sky130_fd_sc_hd__or4_2
X_4379_ VGND VPWR VPWR VGND _3878_ _3876_ _3857_ _3917_ ZI_sky130_fd_sc_hd__or3_2
X_7167_ VGND VPWR VPWR VGND _2615_ _2616_ _2613_ _2617_ ZI_sky130_fd_sc_hd__or3_2
X_7098_ VGND VPWR _2549_ _2546_ _2548_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6118_ VPWR VGND _1580_ _1579_ _1578_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6049_ _1313_ _1511_ _1338_ _1363_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_64_654 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_64_632 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_106_233 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_32_540 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_96_Left_209 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_27_345 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_82_473 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_70_624 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5420_ VGND VPWR VGND VPWR _0889_ _0888_ _0670_ _0613_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_112_225 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5351_ _0546_ _0820_ _0655_ _0645_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8070_ VGND VPWR _3452_ _2323_ _3232_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5282_ VGND VPWR _0648_ _0695_ _0752_ _0751_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
X_4302_ VGND VPWR VGND VPWR _3840_ new_block[38] sword_ctr_reg\[1\] sword_ctr_reg\[0\]
+ ZI_sky130_fd_sc_hd__and3b_2
X_7021_ VPWR VGND VPWR VGND _2285_ _2260_ _2097_ _2208_ _2473_ ZI_sky130_fd_sc_hd__a22o_2
X_4233_ VGND VPWR _3776_ _3775_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7923_ VPWR VGND VPWR VGND _3309_ _3257_ _3318_ _3237_ _0992_ _3319_ ZI_sky130_fd_sc_hd__a221o_2
X_7854_ VGND VPWR _3257_ _0161_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_81_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6805_ VGND VPWR _2259_ _2239_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7785_ VGND VPWR _3194_ _1944_ _3193_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_632 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6736_ VGND VPWR _2190_ _2189_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4997_ VPWR VGND VGND VPWR _0421_ _0466_ _0467_ _0468_ _0469_ ZI_sky130_fd_sc_hd__and4b_2
XFILLER_0_33_337 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_45_197 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6667_ VGND VPWR VGND VPWR _2059_ _2054_ _3832_ _2121_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_60_123 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6598_ VGND VPWR VGND VPWR _2052_ sword_ctr_reg\[0\] new_block[93] sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__and3b_2
X_8406_ VGND VPWR VPWR VGND clk _0008_ reset_n round[1] ZI_sky130_fd_sc_hd__dfrtp_2
X_5618_ VPWR VGND VPWR VGND _0846_ _0731_ _0666_ _0661_ _1084_ ZI_sky130_fd_sc_hd__a22o_2
X_5549_ VGND VPWR VPWR VGND _1014_ _1015_ _0693_ _1016_ ZI_sky130_fd_sc_hd__or3_2
X_8337_ VPWR VGND VPWR VGND _3694_ round_key[25] block[25] ZI_sky130_fd_sc_hd__or2_2
X_8268_ VPWR VGND _3631_ _0904_ _0809_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8199_ VGND VPWR _3569_ _3566_ _3568_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7219_ VPWR VGND VPWR VGND _2665_ _2667_ _2666_ _2664_ _2668_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_28_109 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_107_553 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_91_281 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_52_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_101_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_107_597 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4920_ VPWR VGND VGND VPWR _0393_ _4008_ _3900_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_59_245 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4851_ VGND VPWR VGND VPWR _3816_ _3933_ _4116_ _4110_ _0325_ ZI_sky130_fd_sc_hd__o22a_2
XFILLER_0_7_548 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7570_ VGND VPWR VGND VPWR _2997_ new_block[82] _2996_ _2993_ _1750_ _0061_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_27_142 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_51_87 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4782_ VGND VPWR VGND VPWR _0256_ _4154_ _0257_ _3949_ ZI_sky130_fd_sc_hd__a21oi_2
X_6521_ VPWR VGND VPWR VGND _1875_ _1877_ _1876_ _1805_ _1977_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_43_624 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_15_337 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6452_ VPWR VGND VPWR VGND _1281_ _1909_ _1908_ _0816_ _1907_ _1910_ ZI_sky130_fd_sc_hd__a221o_2
X_5403_ VPWR VGND VPWR VGND _0825_ _0748_ _0606_ _0692_ _0872_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_2_253 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6383_ VPWR VGND VPWR VGND _1281_ _0524_ _1841_ _0816_ _1840_ _1842_ ZI_sky130_fd_sc_hd__a221o_2
X_8122_ VPWR VGND _3500_ block[100] round_key[100] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_2_297 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5334_ VGND VPWR _0804_ _0798_ _0803_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8053_ VGND VPWR _3437_ _0907_ _1058_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5265_ VPWR VGND VPWR VGND _0735_ _0734_ ZI_sky130_fd_sc_hd__inv_2
X_5196_ VGND VPWR _0666_ _0665_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7004_ _2199_ _2456_ _2252_ _2175_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_4216_ VPWR VGND VPWR VGND _3762_ sword_ctr_reg\[0\] ZI_sky130_fd_sc_hd__inv_2
X_7906_ VPWR VGND _3303_ _0241_ _0480_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7837_ VGND VPWR _3241_ _2416_ _2497_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_38_407 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7768_ VPWR VGND VPWR VGND _3150_ _3159_ _3178_ _3139_ _1057_ _3179_ ZI_sky130_fd_sc_hd__a221o_2
X_7699_ VGND VPWR _3116_ _4069_ _0306_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6719_ VPWR VGND VGND VPWR _2110_ _2173_ _2128_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_34_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_33_178 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_104_545 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_104_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_112_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_24_112 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_21_57 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_97_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5050_ VGND VPWR VPWR VGND _0519_ _0516_ _0521_ _0444_ _0520_ ZI_sky130_fd_sc_hd__o211a_2
X_5952_ VGND VPWR _1414_ _1413_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4903_ VPWR VGND _0377_ _0376_ _4076_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5883_ VPWR VGND VGND VPWR _1344_ _1345_ _1307_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_75_546 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_7_301 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7622_ VGND VPWR _3045_ _1908_ _2691_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4834_ VGND VPWR _0309_ _0149_ _0308_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7553_ VGND VPWR VGND VPWR _2981_ _2980_ _2982_ _2642_ ZI_sky130_fd_sc_hd__a21oi_2
X_4765_ VPWR VGND _0241_ round_key[65] new_block[65] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_7_389 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_16_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6504_ VPWR VGND _1961_ new_block[117] round_key[117] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_15_156 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_43_465 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7484_ VGND VPWR _2919_ _1681_ _1825_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4696_ VGND VPWR VGND VPWR _0171_ _3949_ _4131_ _3918_ _0172_ ZI_sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_30_137 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6435_ VGND VPWR _1893_ _1890_ _1892_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6366_ VGND VPWR _1825_ _1576_ _1762_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8105_ VGND VPWR _3484_ _2410_ _2551_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5317_ VGND VPWR _0787_ _0677_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8036_ VGND VPWR VGND VPWR _3419_ _0444_ _3421_ _3422_ ZI_sky130_fd_sc_hd__a21o_2
X_6297_ VGND VPWR _1757_ _1577_ _1756_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5248_ VPWR VGND _0616_ _0718_ _0717_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5179_ VGND VPWR VGND VPWR _0543_ _0537_ _0649_ _3880_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_66_502 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_66_524 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_21_126 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_107_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_72_527 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_25_432 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_25_443 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_37_281 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_106_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4550_ VPWR VGND VPWR VGND dec_ctrl_reg\[2\] _3759_ _3766_ dec_ctrl_reg\[1\] _4088_
+ ZI_sky130_fd_sc_hd__or4_2
X_4481_ VPWR VGND VGND VPWR _3803_ _4019_ _3851_ ZI_sky130_fd_sc_hd__nor2_2
X_6220_ VGND VPWR _1681_ _1679_ _1680_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6151_ VPWR VGND VPWR VGND _1607_ _1611_ _1612_ _1599_ _1601_ ZI_sky130_fd_sc_hd__or4b_2
X_5102_ VGND VPWR VGND VPWR new_block[8] sword_ctr_reg\[0\] _0572_ sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__nand3_2
X_6082_ VPWR VGND VGND VPWR _1524_ _1544_ _1507_ ZI_sky130_fd_sc_hd__nor2_2
X_5033_ VGND VPWR VGND VPWR _4131_ _3906_ _0504_ _3882_ ZI_sky130_fd_sc_hd__a21oi_2
X_6984_ VGND VPWR VGND VPWR _2435_ _2186_ _2126_ _2157_ _2436_ ZI_sky130_fd_sc_hd__a31o_2
X_5935_ VGND VPWR _1397_ _1396_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5866_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[116] sword_ctr_reg\[0\] _1328_
+ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_63_505 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7605_ VGND VPWR VGND VPWR _3030_ _3029_ _3027_ _3025_ ZI_sky130_fd_sc_hd__o21a_2
X_4817_ VGND VPWR VGND VPWR _0292_ _0291_ _0288_ _0285_ _3958_ ZI_sky130_fd_sc_hd__and4_2
XFILLER_0_90_302 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_7_153 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_28_292 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5797_ VPWR VGND VPWR VGND _1035_ _1159_ _1092_ _1034_ _1260_ ZI_sky130_fd_sc_hd__or4_2
X_7536_ VGND VPWR VGND VPWR _2967_ _2966_ _2965_ _2963_ ZI_sky130_fd_sc_hd__o21a_2
X_4748_ VGND VPWR VGND VPWR _3925_ _3945_ _4138_ _4135_ _0224_ _3919_ ZI_sky130_fd_sc_hd__a2111o_2
X_4679_ VGND VPWR _0156_ _0152_ _0155_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7467_ VPWR VGND _2903_ _2883_ _1763_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_1_Right_1 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6418_ VPWR VGND VPWR VGND _1408_ _1493_ _1359_ _1433_ _1876_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_101_301 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7398_ VGND VPWR _2840_ _2837_ _2839_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6349_ VPWR VGND VGND VPWR _1372_ _1519_ _1515_ _1474_ _1440_ _1808_ ZI_sky130_fd_sc_hd__a311o_2
X_8019_ VGND VPWR _3406_ _2788_ _3405_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_343 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_54_527 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_19_281 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_10_608 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_94_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_630 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_76_129 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5720_ VGND VPWR _1185_ _1138_ _1184_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_332 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_45_505 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5651_ VPWR VGND VPWR VGND _0722_ _0834_ _0740_ _0692_ _1117_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_4_123 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8370_ VPWR VGND _3723_ _1578_ _1569_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4602_ VGND VPWR VGND VPWR _4139_ _3949_ _4138_ _3873_ ZI_sky130_fd_sc_hd__o21a_2
X_5582_ VPWR VGND VGND VPWR _0723_ _1049_ _0774_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_25_273 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_53_593 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7321_ VPWR VGND VPWR VGND _2115_ _2279_ _2123_ _2154_ _2768_ ZI_sky130_fd_sc_hd__a22o_2
X_4533_ VGND VPWR _4071_ _4065_ _4070_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7252_ VGND VPWR VPWR VGND _2699_ _2688_ _2701_ _1277_ _2700_ ZI_sky130_fd_sc_hd__o211a_2
X_6203_ VPWR VGND VPWR VGND _1661_ _1663_ _1662_ _1660_ _1664_ ZI_sky130_fd_sc_hd__or4_2
X_4464_ _3803_ _4002_ _3857_ _3869_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_68_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7183_ VGND VPWR _2633_ _2309_ _2560_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4395_ VGND VPWR _3933_ _3887_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6134_ VGND VPWR VGND VPWR _1464_ _1522_ _1592_ _1593_ _1595_ _1594_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_110_197 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6065_ VPWR VGND VGND VPWR _1357_ _1527_ _1344_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_30_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5016_ VPWR VGND _0488_ block[70] round_key[70] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6967_ VPWR VGND _2420_ block[121] round_key[121] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5918_ _1300_ _1380_ _3752_ _1305_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_48_365 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6898_ VPWR VGND VPWR VGND _2337_ _2350_ _2342_ _2271_ _2351_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_75_162 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5849_ VGND VPWR VGND VPWR new_block[87] _3763_ _3797_ _1309_ _1311_ _1310_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_48_398 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_90_132 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_63_346 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_106_448 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_91_666 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_90_165 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7519_ VGND VPWR _2951_ _1900_ _2950_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8499_ VGND VPWR VPWR VGND clk _0101_ reset_n new_block[58] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_31_254 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_12_490 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_39_376 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_10_416 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7870_ VGND VPWR _3271_ _1055_ _2987_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6821_ VPWR VGND _2141_ _2275_ _2235_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_9_215 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_58_641 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_9_237 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6752_ VGND VPWR VGND VPWR _2206_ _2204_ _2203_ _2205_ _2158_ _2188_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_73_600 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_70_42 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5703_ VGND VPWR VGND VPWR _1168_ _0841_ _0722_ _0666_ _0701_ _0754_ ZI_sky130_fd_sc_hd__a32o_2
X_6683_ VGND VPWR VGND VPWR _2137_ _2132_ _2127_ _2107_ _2136_ _2073_ ZI_sky130_fd_sc_hd__a32o_2
X_8422_ VGND VPWR VPWR VGND clk _0024_ reset_n new_block[109] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_70_97 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5634_ VGND VPWR VGND VPWR _1100_ _0571_ _0580_ _0619_ _0841_ _0674_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_5_432 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8353_ VGND VPWR _3708_ _3706_ _3707_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_243 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5565_ VPWR VGND VPWR VGND _0844_ _1031_ _0947_ _0892_ _1032_ ZI_sky130_fd_sc_hd__or4_2
X_7304_ VGND VPWR VGND VPWR _2361_ _2343_ _2288_ _2681_ _2751_ _2750_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_78_3 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8284_ VPWR VGND _3646_ _3418_ _0987_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4516_ VPWR VGND VGND VPWR _3941_ _3921_ _4054_ _3917_ _3961_ ZI_sky130_fd_sc_hd__o22ai_2
X_5496_ VPWR VGND _0846_ _0964_ _0763_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_7235_ VPWR VGND VPWR VGND _2681_ _2683_ _2682_ _2680_ _2684_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_111_462 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4447_ VPWR VGND VGND VPWR _3984_ _3985_ _3982_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_0_181 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_111_495 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7166_ VPWR VGND VPWR VGND _2234_ _2246_ _2155_ _2233_ _2236_ _2616_ ZI_sky130_fd_sc_hd__a221o_2
X_6117_ VPWR VGND _1579_ round_key[8] new_block[8] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4378_ VGND VPWR VPWR VGND _3891_ _3915_ _3890_ _3916_ ZI_sky130_fd_sc_hd__or3_2
X_7097_ VPWR VGND _2548_ _2547_ _2316_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6048_ VPWR VGND VGND VPWR _1307_ _1510_ _1288_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_95_202 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7999_ VGND VPWR _3388_ _3386_ _3387_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_666 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_44_390 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_106_289 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_40_23 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_55_666 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_54_187 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5350_ VGND VPWR VGND VPWR _4104_ new_block[104] _0819_ _0815_ _0793_ _0019_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_112_237 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_10_235 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5281_ VPWR VGND _0579_ _0751_ _0639_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_4301_ sword_ctr_reg\[1\] _3839_ sword_ctr_reg\[0\] new_block[6] VPWR VGND VPWR VGND
+ ZI_sky130_fd_sc_hd__and3_2
X_7020_ VPWR VGND VPWR VGND _2208_ _2279_ _2144_ _2255_ _2472_ ZI_sky130_fd_sc_hd__a22o_2
X_4232_ VGND VPWR _3775_ _3774_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_4_67 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_65_75 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7922_ VPWR VGND _3318_ block[82] round_key[82] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7853_ VPWR VGND _3256_ block[107] round_key[107] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6804_ VGND VPWR VGND VPWR _2258_ _2171_ _2230_ _2254_ _2257_ ZI_sky130_fd_sc_hd__a211o_2
X_7784_ VGND VPWR _3193_ _1571_ _1764_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4996_ VGND VPWR VGND VPWR _3862_ _3992_ _3990_ _4153_ _0468_ ZI_sky130_fd_sc_hd__o22a_2
XFILLER_0_14_90 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_105_81 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6735_ VPWR VGND VGND VPWR _2095_ _2189_ _2188_ ZI_sky130_fd_sc_hd__nor2_2
X_6666_ VGND VPWR _2120_ _2119_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8405_ VGND VPWR VPWR VGND clk _0007_ reset_n round[0] ZI_sky130_fd_sc_hd__dfrtp_2
X_6597_ VGND VPWR VGND VPWR _2051_ new_block[61] sword_ctr_reg\[1\] sword_ctr_reg\[0\]
+ ZI_sky130_fd_sc_hd__and3b_2
X_5617_ VGND VPWR VGND VPWR _0636_ _0923_ _1079_ _1080_ _1083_ _1082_ ZI_sky130_fd_sc_hd__a2111o_2
X_5548_ VGND VPWR VGND VPWR _1015_ _0713_ _0728_ _0975_ ZI_sky130_fd_sc_hd__o21a_2
X_8336_ VPWR VGND VGND VPWR _3693_ round_key[25] block[25] ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_60_168 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8267_ VGND VPWR _3630_ _0909_ _1059_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_393 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5479_ VGND VPWR VGND VPWR _0947_ _0851_ _0644_ _0606_ _0612_ _0704_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_111_281 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7218_ _2265_ _2667_ _2188_ _2212_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8198_ VGND VPWR _3568_ _3334_ _3567_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7149_ VPWR VGND VPWR VGND _2150_ _2223_ _2599_ _2336_ _2158_ ZI_sky130_fd_sc_hd__a22oi_2
XFILLER_0_49_482 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_36_121 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_64_430 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_10_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_101_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_20_599 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4850_ VPWR VGND VPWR VGND _4130_ _0323_ _4146_ _0322_ _0324_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_59_257 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_28_622 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_51_22 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6520_ VPWR VGND VPWR VGND _1481_ _1975_ _1482_ _1476_ _1976_ ZI_sky130_fd_sc_hd__or4_2
X_4781_ VPWR VGND VGND VPWR _0256_ _3934_ _3925_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_82_293 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6451_ VGND VPWR _1909_ _0168_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6382_ VPWR VGND _1841_ new_block[115] round_key[115] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5402_ VGND VPWR VGND VPWR _0871_ _0734_ _0656_ _0635_ _0664_ _0580_ ZI_sky130_fd_sc_hd__a32o_2
X_5333_ VGND VPWR _0803_ _0799_ _0802_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8121_ VPWR VGND VGND VPWR _3498_ _3499_ _3497_ ZI_sky130_fd_sc_hd__nor2_2
X_8052_ VPWR VGND _3436_ _3414_ _2849_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5264_ VPWR VGND VGND VPWR _0595_ _0734_ _0620_ ZI_sky130_fd_sc_hd__nor2_2
X_5195_ VPWR VGND _0544_ _0665_ _0638_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_7003_ VGND VPWR VGND VPWR _2455_ _2345_ _2265_ _2285_ ZI_sky130_fd_sc_hd__o21a_2
X_4215_ VPWR VGND VPWR VGND _3761_ next ZI_sky130_fd_sc_hd__inv_2
XFILLER_0_76_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7905_ VGND VPWR VGND VPWR _3240_ new_block[48] _3302_ _3300_ _1562_ _0091_ ZI_sky130_fd_sc_hd__o32a_2
X_7836_ VGND VPWR VGND VPWR _3240_ new_block[41] _3239_ _3236_ _0899_ _0084_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_19_600 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7767_ VPWR VGND _3178_ block[3] round_key[3] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4979_ VPWR VGND VPWR VGND _4042_ _4031_ _3898_ _3938_ _0451_ ZI_sky130_fd_sc_hd__a22o_2
X_7698_ VGND VPWR _3115_ _3110_ _3114_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6718_ VPWR VGND VPWR VGND _2158_ _2171_ _2102_ _2169_ _2172_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_61_411 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_6_560 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_18_187 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_33_113 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6649_ VPWR VGND VGND VPWR _3880_ _2089_ _2094_ _2103_ ZI_sky130_fd_sc_hd__nor3_2
XFILLER_0_14_360 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_104_557 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8319_ VPWR VGND VGND VPWR _1568_ _3678_ _4089_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_71_208 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_64_282 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_40_606 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_46_22 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5951_ VGND VPWR VGND VPWR _1329_ _1324_ _3832_ _1413_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_99_190 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4902_ VPWR VGND _0376_ round_key[76] new_block[76] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5882_ VGND VPWR _1344_ _1343_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_47_238 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4833_ VPWR VGND _0308_ round_key[83] new_block[83] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7621_ VPWR VGND _3044_ _3043_ _1241_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7552_ VGND VPWR _2981_ _2316_ _2557_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4764_ VGND VPWR _0240_ _0142_ _0239_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6503_ VPWR VGND _1960_ block[21] round_key[21] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7483_ VGND VPWR _2918_ _2913_ _2917_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_477 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6434_ VGND VPWR _1892_ _1568_ _1891_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4695_ VPWR VGND VPWR VGND _0171_ _4148_ _4190_ ZI_sky130_fd_sc_hd__or2_2
XFILLER_0_31_639 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6365_ VGND VPWR _1824_ _1577_ _1755_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_87_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8104_ VGND VPWR _3483_ _2999_ _3482_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5316_ VPWR VGND _0785_ _0786_ _0741_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_6296_ VPWR VGND _1756_ _1755_ _1689_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5247_ VGND VPWR _0717_ _0716_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8035_ VPWR VGND VPWR VGND _3149_ _4093_ _3420_ _2702_ _1137_ _3421_ ZI_sky130_fd_sc_hd__a221o_2
X_5178_ VGND VPWR _0648_ _0644_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7819_ VPWR VGND _3225_ _3224_ _3223_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_108_137 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_34_411 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_34_477 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_104_321 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_107_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_89_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_69_385 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_13_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_12_105 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_12_116 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4480_ VGND VPWR VGND VPWR _4013_ _4012_ _4014_ _4015_ _4018_ _4017_ ZI_sky130_fd_sc_hd__a2111o_2
X_6150_ VPWR VGND VGND VPWR _1460_ _1384_ _1507_ _1547_ _1611_ _1610_ ZI_sky130_fd_sc_hd__o221a_2
XFILLER_0_20_171 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5101_ VGND VPWR _0571_ _0570_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6081_ VPWR VGND VGND VPWR _1479_ _1543_ _1447_ ZI_sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_29_Left_142 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5032_ VGND VPWR VGND VPWR _4023_ _3816_ _0503_ _3955_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_57_98 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_79_105 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6983_ _2182_ _2435_ _2252_ _2199_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5934_ _1318_ _1396_ _1312_ _1377_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5865_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] _1327_ new_block[84] ZI_sky130_fd_sc_hd__and2b_2
XPHY_EDGE_ROW_38_Left_151 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_7_121 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7604_ VGND VPWR VGND VPWR _3027_ _3025_ _3029_ _3028_ ZI_sky130_fd_sc_hd__a21oi_2
X_4816_ VPWR VGND VPWR VGND _0291_ _3877_ _3976_ _3910_ _0289_ _0290_ ZI_sky130_fd_sc_hd__o311a_2
X_5796_ VPWR VGND VPWR VGND _1247_ _1258_ _1255_ _1203_ _1259_ ZI_sky130_fd_sc_hd__or4_2
X_7535_ VGND VPWR VGND VPWR _2965_ _2963_ _2966_ _2642_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_71_561 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4747_ VPWR VGND VPWR VGND _4056_ _0222_ _0223_ _3866_ _4049_ ZI_sky130_fd_sc_hd__or4b_2
XFILLER_0_31_436 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7466_ VGND VPWR VGND VPWR _2894_ new_block[73] _2902_ _2900_ _0899_ _0052_ ZI_sky130_fd_sc_hd__o32a_2
X_4678_ VPWR VGND _0155_ _0154_ _0153_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_3_360 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7397_ VGND VPWR _2839_ _1127_ _2838_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6417_ VGND VPWR VGND VPWR _1487_ _1538_ _1875_ _1384_ ZI_sky130_fd_sc_hd__a21oi_2
X_6348_ VPWR VGND VPWR VGND _1641_ _1806_ _1803_ _1457_ _1807_ ZI_sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_47_Left_160 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6279_ VPWR VGND VGND VPWR _1739_ _1736_ _1738_ ZI_sky130_fd_sc_hd__nand2_2
X_8018_ VPWR VGND _3405_ _2845_ _0810_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_39_525 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_105_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_85_642 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5650_ VGND VPWR VGND VPWR _1116_ _0656_ _0825_ _0763_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_45_517 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_84_141 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_38_580 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4601_ VPWR VGND VGND VPWR _3962_ _4138_ _4115_ ZI_sky130_fd_sc_hd__nor2_2
X_5581_ VGND VPWR VGND VPWR _1048_ _0775_ _0689_ _1046_ _1047_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_4_135 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_13_403 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7320_ VPWR VGND VPWR VGND _2766_ _2187_ _2230_ _2107_ _2233_ _2767_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_108_490 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4532_ VGND VPWR _4070_ _4066_ _4069_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7251_ VPWR VGND VGND VPWR _2700_ _2688_ _2699_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_111_600 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4463_ VGND VPWR VGND VPWR _3903_ _3997_ _4000_ _4001_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_7_67 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6202_ VGND VPWR VGND VPWR _1663_ _1443_ _1434_ _1360_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_68_53 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_15_Right_15 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7182_ VGND VPWR _2632_ _2310_ _2487_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4394_ VGND VPWR _3932_ _3860_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6133_ VPWR VGND _1452_ _1594_ _1528_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_6064_ VGND VPWR VGND VPWR _1525_ _1521_ _1522_ _1523_ _1526_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_84_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5015_ VGND VPWR VPWR VGND _0485_ _0484_ _0487_ _0444_ _0486_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_23_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_84_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6966_ VGND VPWR VPWR VGND _2417_ _2415_ _2419_ _1277_ _2418_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_76_620 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5917_ VGND VPWR _1379_ _1378_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_75_130 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_48_355 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6897_ VPWR VGND VGND VPWR _2349_ _2348_ _2118_ _2199_ _2233_ _2350_ ZI_sky130_fd_sc_hd__a311o_2
X_5848_ sword_ctr_reg\[1\] _1310_ sword_ctr_reg\[0\] new_block[23] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
X_5779_ VGND VPWR VGND VPWR _1009_ new_block[110] _1242_ _1239_ _1227_ _0025_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_44_572 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7518_ VGND VPWR _2950_ _1578_ _1819_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8498_ VGND VPWR VPWR VGND clk _0100_ reset_n new_block[57] ZI_sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_33_Right_33 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_101_121 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7449_ VGND VPWR _2887_ _1683_ _1832_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_42_Right_42 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_39_311 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_109_221 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_66_141 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_82_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Right_60 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_89_244 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6820_ VGND VPWR VGND VPWR _2274_ _2169_ _2273_ _2135_ _2215_ _2252_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_9_249 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6751_ VPWR VGND VGND VPWR _2146_ _2205_ _2128_ ZI_sky130_fd_sc_hd__nor2_2
X_5702_ VPWR VGND VPWR VGND _1044_ _1166_ _1163_ _0882_ _1167_ ZI_sky130_fd_sc_hd__or4_2
X_6682_ VGND VPWR _2136_ _2135_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8421_ VGND VPWR VPWR VGND clk _0023_ reset_n new_block[108] ZI_sky130_fd_sc_hd__dfrtp_2
X_5633_ VGND VPWR VGND VPWR _0787_ _0651_ _0685_ _0833_ _1099_ _0653_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_5_444 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5564_ VPWR VGND VPWR VGND _1031_ _1029_ _1030_ ZI_sky130_fd_sc_hd__or2_2
X_8352_ VPWR VGND _3707_ _1764_ _1677_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_72_166 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_5_488 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4515_ VGND VPWR VPWR VGND _3849_ _4053_ _3917_ _4052_ _4022_ ZI_sky130_fd_sc_hd__a31oi_2
X_7303_ VPWR VGND VPWR VGND _2294_ _2107_ _2259_ _2327_ _2256_ _2750_ ZI_sky130_fd_sc_hd__a221o_2
X_8283_ VGND VPWR _3645_ _3642_ _3644_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_553 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_103_Right_103 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5495_ VPWR VGND VGND VPWR _0652_ _0963_ _0856_ ZI_sky130_fd_sc_hd__nor2_2
X_7234_ VGND VPWR VGND VPWR _2299_ _2297_ _2271_ _2269_ _2683_ _2116_ ZI_sky130_fd_sc_hd__a2111o_2
X_4446_ VGND VPWR _3984_ _3983_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_111_474 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7165_ VGND VPWR VGND VPWR _2615_ _2202_ _2233_ _2363_ _2614_ ZI_sky130_fd_sc_hd__a211o_2
X_4377_ VGND VPWR VGND VPWR _3915_ _3843_ _3884_ _3883_ _3914_ ZI_sky130_fd_sc_hd__o211ai_2
XFILLER_0_0_193 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_95_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6116_ VPWR VGND _1578_ round_key[13] new_block[13] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7096_ VPWR VGND _2547_ _2048_ _1841_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6047_ VGND VPWR VGND VPWR _1509_ _1443_ _1419_ _1506_ _1508_ ZI_sky130_fd_sc_hd__a211o_2
X_7998_ VPWR VGND _3387_ _0997_ _0807_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_95_225 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6949_ VPWR VGND VPWR VGND _2399_ _2401_ _2400_ _2398_ _2402_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_64_612 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_17_561 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_106_246 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_54_100 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_112_249 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5280_ VPWR VGND VPWR VGND _0749_ _0607_ _0710_ _0747_ _0748_ _0750_ ZI_sky130_fd_sc_hd__a221o_2
X_4300_ VGND VPWR _3838_ _3837_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_10_247 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4231_ VGND VPWR _3774_ _3773_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_4_79 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_65_43 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7921_ VGND VPWR VPWR VGND _3315_ _3314_ _3317_ _3265_ _3316_ ZI_sky130_fd_sc_hd__o211a_2
X_7852_ VGND VPWR VPWR VGND _3253_ _3252_ _3255_ _3118_ _3254_ ZI_sky130_fd_sc_hd__o211a_2
X_6803_ VPWR VGND VPWR VGND _2256_ _2255_ _2115_ _2143_ _2257_ ZI_sky130_fd_sc_hd__a22o_2
X_7783_ VPWR VGND _3192_ _3191_ _1757_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_58_450 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4995_ VGND VPWR VGND VPWR _3930_ _3874_ _3993_ _4140_ _0467_ ZI_sky130_fd_sc_hd__o22a_2
X_6734_ VPWR VGND VGND VPWR _2188_ _3754_ _2160_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_18_336 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_45_122 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_46_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_90_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6665_ VPWR VGND VGND VPWR _2110_ _2119_ _2118_ ZI_sky130_fd_sc_hd__nor2_2
X_8404_ VGND VPWR VPWR VGND clk _0006_ reset_n sword_ctr_reg\[1\] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_520 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5616_ VPWR VGND VPWR VGND _0863_ _1081_ _0820_ _0715_ _1082_ ZI_sky130_fd_sc_hd__or4_2
X_6596_ sword_ctr_reg\[1\] _2050_ sword_ctr_reg\[0\] new_block[29] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
X_5547_ VGND VPWR VGND VPWR _1014_ _0763_ _0583_ _0606_ _0767_ _0886_ ZI_sky130_fd_sc_hd__a32o_2
X_8335_ VGND VPWR VPWR VGND _3690_ _1896_ _3692_ _0366_ _3691_ ZI_sky130_fd_sc_hd__o211a_2
X_8266_ VGND VPWR VGND VPWR _3548_ new_block[18] _3629_ _3627_ _1750_ _0125_ ZI_sky130_fd_sc_hd__o32a_2
X_5478_ VPWR VGND VPWR VGND _0615_ _0692_ _0785_ _0670_ _0946_ ZI_sky130_fd_sc_hd__a22o_2
X_7217_ VGND VPWR VGND VPWR _2666_ _2106_ _2177_ _2184_ ZI_sky130_fd_sc_hd__o21a_2
X_4429_ VPWR VGND VGND VPWR _3967_ _3948_ _3804_ ZI_sky130_fd_sc_hd__nand2_2
X_8197_ VGND VPWR _3567_ _0240_ _0312_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7148_ VPWR VGND VPWR VGND _2120_ _2246_ _2299_ _2372_ _2598_ ZI_sky130_fd_sc_hd__a22o_2
X_7079_ VPWR VGND VPWR VGND _2520_ _2529_ _2524_ _2365_ _2530_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_96_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_36_133 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_51_169 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_19_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_51_34 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_74_228 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4780_ VPWR VGND VPWR VGND _0254_ _4189_ _4019_ _4010_ _3934_ _0255_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_55_431 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_82_272 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_70_412 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6450_ VPWR VGND _1908_ new_block[116] round_key[116] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_43_659 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6381_ VPWR VGND _1840_ block[19] round_key[19] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5401_ VGND VPWR VGND VPWR _0851_ _0645_ _0778_ _0870_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_30_309 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5332_ VGND VPWR _0802_ _0800_ _0801_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8120_ VGND VPWR VGND VPWR _3496_ _3495_ _0158_ _3498_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_2_277 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Left_123 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8051_ VGND VPWR VGND VPWR _3150_ _4094_ _3433_ _3434_ _3435_ ZI_sky130_fd_sc_hd__a31o_2
X_5263_ VGND VPWR VPWR VGND _0730_ _0732_ _0725_ _0733_ ZI_sky130_fd_sc_hd__or3_2
X_5194_ VGND VPWR _0664_ _0663_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7002_ VGND VPWR VGND VPWR _2454_ _2373_ _2205_ _2120_ ZI_sky130_fd_sc_hd__o21a_2
X_4214_ VGND VPWR VGND VPWR _0003_ _3758_ _3756_ _3760_ dec_ctrl_reg\[2\] ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_92_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7904_ VPWR VGND VPWR VGND _3219_ _3257_ _3301_ _3237_ _0809_ _3302_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_92_85 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7835_ VGND VPWR _3240_ _3152_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_19_612 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_65_228 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7766_ VPWR VGND VGND VPWR _3176_ _3177_ _3175_ ZI_sky130_fd_sc_hd__nor2_2
X_4978_ VGND VPWR VGND VPWR _0450_ _4008_ _4148_ _0449_ ZI_sky130_fd_sc_hd__o21a_2
X_7697_ VPWR VGND _3114_ _3113_ _0382_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6717_ VGND VPWR _2171_ _2170_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_33_136 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_104_503 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6648_ VGND VPWR _2102_ _2101_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6579_ VPWR VGND VGND VPWR _1466_ _2034_ _1445_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_104_569 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8318_ VPWR VGND VPWR VGND _3677_ round_key[55] block[55] ZI_sky130_fd_sc_hd__or2_2
X_8249_ VGND VPWR _3614_ _1062_ _3613_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_25_604 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_52_412 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_12_309 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_52_489 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_46_34 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5950_ VPWR VGND VGND VPWR _1412_ _1368_ _1381_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_1_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4901_ VGND VPWR _0375_ _0373_ _0374_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5881_ VGND VPWR VPWR VGND _1287_ _1294_ _3879_ _1343_ ZI_sky130_fd_sc_hd__or3_2
X_7620_ VPWR VGND _3043_ _1280_ _1146_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_87_386 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_62_66 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4832_ VGND VPWR _0307_ _4075_ _4072_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7551_ VGND VPWR _2980_ _2978_ _2979_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4763_ VGND VPWR _0239_ _4061_ _0238_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_261 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6502_ VGND VPWR _1959_ _0161_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_83_581 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7482_ VGND VPWR _2917_ _2914_ _2916_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4694_ VGND VPWR VGND VPWR _4104_ new_block[97] _0170_ _0160_ _0140_ _0012_ ZI_sky130_fd_sc_hd__o32a_2
X_6433_ VPWR VGND _1891_ round_key[19] new_block[19] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_11_70 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_43_489 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_101_539 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6364_ VGND VPWR _1823_ _1818_ _1822_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8103_ VPWR VGND _3482_ _2560_ _1841_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5315_ VPWR VGND _0581_ _0785_ _0557_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_6295_ VPWR VGND _1755_ round_key[10] new_block[10] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5246_ VPWR VGND VGND VPWR _0655_ _0716_ _0649_ ZI_sky130_fd_sc_hd__nor2_2
X_8034_ VPWR VGND _3420_ block[60] round_key[60] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_89_Right_89 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5177_ VGND VPWR VGND VPWR _0628_ _0546_ _0636_ _0641_ _0647_ _0646_ ZI_sky130_fd_sc_hd__a2111o_2
X_7818_ VPWR VGND _3224_ _2323_ _2309_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_98_Right_98 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_109_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_66_548 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_81_518 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7749_ VPWR VGND _3161_ _1831_ _1820_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_104_300 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_61_242 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_14_191 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_16_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_107_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_89_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_29_206 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_107_160 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_13_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_107_182 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_80_584 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_0_501 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_12_128 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_0_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_20_183 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6080_ VPWR VGND VGND VPWR _1473_ _1542_ _1436_ ZI_sky130_fd_sc_hd__nor2_2
X_5100_ VPWR VGND _0557_ _0570_ _0569_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_110_358 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5031_ VPWR VGND VPWR VGND _0401_ _0469_ _0502_ _0273_ _0348_ ZI_sky130_fd_sc_hd__or4b_2
X_6982_ VGND VPWR VGND VPWR _2171_ _2338_ _2430_ _2431_ _2434_ _2433_ ZI_sky130_fd_sc_hd__a2111o_2
X_5933_ VGND VPWR _1395_ _1394_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_87_161 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5864_ sword_ctr_reg\[1\] _1326_ sword_ctr_reg\[0\] new_block[20] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_8_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4815_ VGND VPWR VGND VPWR _3862_ _3896_ _4114_ _3969_ _0290_ ZI_sky130_fd_sc_hd__o22a_2
X_7603_ VGND VPWR _3028_ _4085_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7534_ VGND VPWR _2965_ _2040_ _2964_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5795_ VGND VPWR VPWR VGND _1256_ _1257_ _0840_ _1258_ ZI_sky130_fd_sc_hd__or3_2
X_4746_ VGND VPWR VGND VPWR _3905_ _3859_ _4036_ _3930_ _3948_ _0222_ ZI_sky130_fd_sc_hd__o32a_2
X_4677_ VPWR VGND _0154_ round_key[73] new_block[73] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7465_ VPWR VGND VPWR VGND _2892_ _2786_ _2901_ _2880_ _0154_ _2902_ ZI_sky130_fd_sc_hd__a221o_2
X_7396_ VPWR VGND _2838_ _2801_ _1188_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_12_640 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6416_ VGND VPWR VGND VPWR _1866_ _1874_ _1870_ _1873_ _1868_ ZI_sky130_fd_sc_hd__and4bb_2
X_6347_ VGND VPWR VGND VPWR _1361_ _1351_ _1698_ _1804_ _1806_ _1805_ ZI_sky130_fd_sc_hd__a2111o_2
X_6278_ VGND VPWR VPWR VGND _1738_ _1390_ _1384_ _1401_ _1737_ ZI_sky130_fd_sc_hd__o31a_2
X_8017_ VGND VPWR _3404_ _1062_ _1138_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5229_ _0591_ _0699_ _0698_ _0626_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_81_337 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_22_415 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_34_253 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_105_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_104_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_104_152 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_30_470 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_43_35 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_85_654 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_84_153 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_45_529 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_84_197 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4600_ VPWR VGND VPWR VGND _4132_ _4136_ _4137_ _4128_ _4130_ ZI_sky130_fd_sc_hd__or4b_2
XFILLER_0_53_540 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5580_ _0571_ _1047_ _0546_ _0735_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_4531_ VPWR VGND _4069_ _4068_ _4067_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7250_ VGND VPWR _2699_ _2690_ _2698_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4462_ VGND VPWR VGND VPWR _3999_ _3998_ _4000_ _3984_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_111_612 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_7_57 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6201_ VGND VPWR VGND VPWR _1399_ _1366_ _1662_ _1487_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_7_79 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7181_ VPWR VGND _2631_ _2630_ _1146_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4393_ VPWR VGND VGND VPWR _3930_ _3931_ _3865_ ZI_sky130_fd_sc_hd__nor2_2
X_6132_ VPWR VGND VGND VPWR _1473_ _1593_ _1538_ ZI_sky130_fd_sc_hd__nor2_2
X_6063_ VPWR VGND VGND VPWR _1524_ _1525_ _1416_ ZI_sky130_fd_sc_hd__nor2_2
X_5014_ VPWR VGND VGND VPWR _0486_ _0484_ _0485_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_84_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6965_ VPWR VGND VGND VPWR _2418_ _2415_ _2417_ ZI_sky130_fd_sc_hd__nand2_2
X_5916_ _1362_ _1378_ _1352_ _1377_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_76_632 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6896_ VGND VPWR VGND VPWR _2349_ _2259_ _2330_ _2168_ _2222_ _2188_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_91_613 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_8_442 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5847_ VGND VPWR VGND VPWR _1309_ new_block[55] sword_ctr_reg\[1\] sword_ctr_reg\[0\]
+ ZI_sky130_fd_sc_hd__and3b_2
X_5778_ VPWR VGND VPWR VGND _4101_ _0524_ _1241_ _0816_ _1240_ _1242_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_106_417 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_16_253 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8497_ VGND VPWR VPWR VGND clk _0099_ reset_n new_block[56] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_44_584 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7517_ VGND VPWR VGND VPWR _2894_ new_block[77] _2949_ _2947_ _1181_ _0056_ ZI_sky130_fd_sc_hd__o32a_2
X_4729_ VPWR VGND VPWR VGND _3997_ _4042_ _4019_ _3925_ _0205_ ZI_sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_2_Left_115 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7448_ VGND VPWR _2886_ _2883_ _2885_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7379_ VPWR VGND _2822_ _1066_ _0914_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_66_120 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_13_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_104_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_82_602 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_66_153 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_54_304 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_81_101 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_66_197 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_109_277 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_82_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_62_392 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_66_Left_179 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_54_34 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6750_ _2100_ _2204_ _2099_ _2182_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5701_ VGND VPWR VGND VPWR _0727_ _0655_ _1090_ _1164_ _1166_ _1165_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_58_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_18_529 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6681_ VGND VPWR _2135_ _2134_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8420_ VGND VPWR VPWR VGND clk _0022_ reset_n new_block[107] ZI_sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_75_Left_188 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5632_ VPWR VGND VPWR VGND _1083_ _1097_ _1089_ _0845_ _1098_ ZI_sky130_fd_sc_hd__or4_2
X_5563_ VPWR VGND VPWR VGND _0739_ _0741_ _0633_ _0701_ _1030_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_41_510 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8351_ VGND VPWR _3706_ _1816_ _1944_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_178 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7302_ VPWR VGND VPWR VGND _2749_ _2716_ _2748_ ZI_sky130_fd_sc_hd__or2_2
X_4514_ VPWR VGND VGND VPWR _4052_ _3898_ _3815_ ZI_sky130_fd_sc_hd__nand2_2
X_8282_ VGND VPWR _3644_ _2838_ _3643_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_267 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5494_ VGND VPWR VGND VPWR _0888_ _0767_ _0958_ _0960_ _0962_ _0961_ ZI_sky130_fd_sc_hd__a2111o_2
X_7233_ VGND VPWR VGND VPWR _2682_ _2202_ _2214_ _2150_ ZI_sky130_fd_sc_hd__o21a_2
X_4445_ VPWR VGND VGND VPWR _3983_ _3869_ _3920_ ZI_sky130_fd_sc_hd__nand2_2
X_4376_ VGND VPWR _3914_ _3752_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7164_ VPWR VGND VPWR VGND _2190_ _2282_ _2136_ _2330_ _2614_ ZI_sky130_fd_sc_hd__a22o_2
X_6115_ VPWR VGND _1577_ round_key[15] new_block[15] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7095_ VPWR VGND _2546_ _2488_ _2312_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_84_Left_197 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6046_ VGND VPWR VGND VPWR _1487_ _1371_ _1508_ _1507_ ZI_sky130_fd_sc_hd__a21oi_2
X_7997_ VGND VPWR _3386_ _3385_ _2825_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_248 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6948_ VPWR VGND VPWR VGND _2138_ _2177_ _2227_ _2195_ _2401_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_48_164 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6879_ VGND VPWR VGND VPWR _2214_ _2330_ _2331_ _2332_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_64_624 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_8_272 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_91_432 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_51_318 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_32_554 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_5_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_99_543 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_24_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_40_47 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_10_215 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_49_67 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4230_ VPWR VGND VGND VPWR _3773_ dec_ctrl_reg\[1\] _3772_ ZI_sky130_fd_sc_hd__nand2_2
X_7920_ VPWR VGND VGND VPWR _3316_ _3314_ _3315_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_65_99 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7851_ VPWR VGND VGND VPWR _3254_ _3252_ _3253_ ZI_sky130_fd_sc_hd__nand2_2
X_6802_ VPWR VGND VGND VPWR _2192_ _2256_ _2146_ ZI_sky130_fd_sc_hd__nor2_2
X_7782_ VGND VPWR _3191_ _3189_ _3190_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4994_ VGND VPWR VGND VPWR _3921_ _3862_ _3961_ _0466_ ZI_sky130_fd_sc_hd__a21o_2
X_6733_ VGND VPWR _2187_ _2186_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_46_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_281 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6664_ VGND VPWR _2118_ _2117_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5615_ VGND VPWR VGND VPWR _0841_ _0859_ _0867_ _1081_ ZI_sky130_fd_sc_hd__a21o_2
X_8403_ VGND VPWR VPWR VGND clk _0005_ reset_n sword_ctr_reg\[0\] ZI_sky130_fd_sc_hd__dfrtp_2
X_6595_ VGND VPWR VGND VPWR _1911_ new_block[119] _2049_ _2046_ _2038_ _0034_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_83_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5546_ VPWR VGND VPWR VGND _1013_ _0940_ _0931_ ZI_sky130_fd_sc_hd__or2_2
X_8334_ VPWR VGND VGND VPWR _3691_ _1896_ _3690_ ZI_sky130_fd_sc_hd__nand2_2
X_8265_ VPWR VGND VPWR VGND _3575_ _3603_ _3628_ _3583_ _1820_ _3629_ ZI_sky130_fd_sc_hd__a221o_2
X_5477_ VPWR VGND VPWR VGND _0942_ _0944_ _0943_ _0941_ _0945_ ZI_sky130_fd_sc_hd__or4_2
X_7216_ VPWR VGND VPWR VGND _2264_ _2176_ _2201_ _2239_ _2665_ ZI_sky130_fd_sc_hd__a22o_2
X_4428_ VPWR VGND VPWR VGND _3838_ _3885_ _3929_ _3831_ _3966_ ZI_sky130_fd_sc_hd__or4_2
X_8196_ VGND VPWR _3566_ _0375_ _3095_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_92_Left_205 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4359_ VPWR VGND VGND VPWR _3896_ _3897_ _3895_ ZI_sky130_fd_sc_hd__nor2_2
X_7147_ VPWR VGND VPWR VGND _2574_ _2596_ _2587_ _2335_ _2597_ ZI_sky130_fd_sc_hd__or4_2
X_7078_ VPWR VGND VGND VPWR _2528_ _2527_ _2127_ _2136_ _2205_ _2529_ ZI_sky130_fd_sc_hd__a311o_2
X_6029_ VPWR VGND VGND VPWR _1490_ _1491_ _1393_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_9_592 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_27_123 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_51_57 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_27_189 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_2_223 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5400_ VGND VPWR VGND VPWR _0648_ _0683_ _0865_ _0866_ _0869_ _0868_ ZI_sky130_fd_sc_hd__a2111o_2
X_6380_ VGND VPWR VGND VPWR _1839_ _1838_ _1837_ _1827_ ZI_sky130_fd_sc_hd__o21a_2
X_5331_ VPWR VGND _0801_ round_key[45] new_block[45] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_2_289 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_11_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8050_ VPWR VGND VPWR VGND _3434_ round_key[62] block[62] ZI_sky130_fd_sc_hd__or2_2
X_5262_ VGND VPWR VGND VPWR _0732_ _0712_ _0612_ _0690_ _0731_ _0688_ ZI_sky130_fd_sc_hd__a32o_2
X_7001_ VGND VPWR VGND VPWR _2171_ _2299_ _2452_ _2133_ _2453_ ZI_sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_76_32 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5193_ VPWR VGND VGND VPWR _0632_ _0663_ _0655_ ZI_sky130_fd_sc_hd__nor2_2
X_4213_ VPWR VGND dec_ctrl_reg\[3\] _3760_ _3759_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_92_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7903_ VPWR VGND _3301_ block[80] round_key[80] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7834_ VPWR VGND VPWR VGND _3219_ _3159_ _3238_ _3237_ _0997_ _3239_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_78_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7765_ VGND VPWR VGND VPWR _3174_ _3170_ _0158_ _3176_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_18_134 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_46_421 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6716_ VPWR VGND _2161_ _2170_ _2129_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_4977_ VPWR VGND VGND VPWR _3978_ _0449_ _3905_ ZI_sky130_fd_sc_hd__nor2_2
X_7696_ VGND VPWR _3113_ _3111_ _3112_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6647_ _2100_ _2101_ _2099_ _2060_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6578_ VPWR VGND VPWR VGND _2030_ _2032_ _2031_ _1637_ _2033_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_33_148 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_104_515 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5529_ VPWR VGND _0997_ round_key[41] new_block[41] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8317_ VPWR VGND VGND VPWR _3676_ round_key[55] block[55] ZI_sky130_fd_sc_hd__nand2_2
X_8248_ VGND VPWR _3613_ _0795_ _0908_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8179_ VPWR VGND _3551_ _0242_ _0238_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_69_579 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_112_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_25_627 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_107_386 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_1_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5880_ VGND VPWR VGND VPWR _1342_ _1332_ _1308_ _1341_ _1337_ _1289_ ZI_sky130_fd_sc_hd__a32o_2
X_4900_ VGND VPWR _0374_ _4074_ _0152_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4831_ VGND VPWR _0306_ _4066_ _0305_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_56 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_7_337 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4762_ VPWR VGND _0238_ round_key[90] new_block[90] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7550_ VGND VPWR _2979_ _0165_ _2632_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_498 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6501_ VGND VPWR VGND VPWR _1958_ _1957_ _1956_ _1954_ ZI_sky130_fd_sc_hd__o21a_2
X_7481_ VGND VPWR _2916_ _1824_ _2915_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4693_ VPWR VGND VPWR VGND _4101_ _0169_ _0165_ _0162_ _0163_ _0170_ ZI_sky130_fd_sc_hd__a221o_2
X_6432_ VGND VPWR _1890_ _1887_ _1889_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_95 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_3_587 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6363_ VGND VPWR _1822_ _1819_ _1821_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8102_ VGND VPWR VGND VPWR _3462_ new_block[2] _3481_ _3479_ _0229_ _0109_ ZI_sky130_fd_sc_hd__o32a_2
X_6294_ VGND VPWR _1754_ _1752_ _1753_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5314_ VPWR VGND VGND VPWR _0783_ _0784_ _0632_ ZI_sky130_fd_sc_hd__nor2_2
X_8033_ VGND VPWR _3419_ _3417_ _3418_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5245_ VPWR VGND _0713_ _0715_ _0709_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5176_ VPWR VGND _0546_ _0646_ _0645_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_19_421 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7817_ VPWR VGND _3223_ _2310_ _1241_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_109_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7748_ VGND VPWR VGND VPWR _3153_ new_block[33] _3160_ _3157_ _0140_ _0076_ ZI_sky130_fd_sc_hd__o32a_2
X_7679_ VPWR VGND _3097_ _3096_ _3095_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_104_378 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_97_630 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_29_218 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_32_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_107_194 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_80_596 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_21_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_40_438 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_57_23 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5030_ VPWR VGND VPWR VGND _0497_ _0500_ _0498_ _0496_ _0501_ ZI_sky130_fd_sc_hd__or4_2
X_6981_ VPWR VGND VPWR VGND _2432_ _2281_ _2143_ _2135_ _2131_ _2433_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_73_33 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5932_ VPWR VGND VGND VPWR _1393_ _1394_ _1391_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_8_602 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5863_ VGND VPWR VGND VPWR _1325_ new_block[52] sword_ctr_reg\[1\] sword_ctr_reg\[0\]
+ ZI_sky130_fd_sc_hd__and3b_2
XFILLER_0_87_184 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4814_ VGND VPWR VGND VPWR _4181_ _4141_ _4023_ _0289_ ZI_sky130_fd_sc_hd__a21o_2
X_5794_ VGND VPWR VPWR VGND _1257_ _0658_ _0696_ _0859_ _0757_ ZI_sky130_fd_sc_hd__o31a_2
X_7602_ VPWR VGND _3027_ _3026_ _0447_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_8_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4745_ VPWR VGND VPWR VGND _0214_ _3908_ _0216_ _0220_ _0221_ ZI_sky130_fd_sc_hd__or4bb_2
X_7533_ VGND VPWR _2964_ _1568_ _1574_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_316 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_71_552 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_98_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4676_ VPWR VGND _0153_ round_key[78] new_block[78] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7464_ VPWR VGND _2901_ block[9] round_key[9] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7395_ VGND VPWR _2837_ _0995_ _2836_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6415_ _1871_ _1873_ _1719_ _1872_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6346_ VPWR VGND VGND VPWR _1445_ _1805_ _1366_ ZI_sky130_fd_sc_hd__nor2_2
X_6277_ VPWR VGND VGND VPWR _1737_ _1527_ _1522_ ZI_sky130_fd_sc_hd__nand2_2
X_8016_ VGND VPWR VGND VPWR _3331_ new_block[58] _3403_ _3401_ _2483_ _0101_ ZI_sky130_fd_sc_hd__o32a_2
X_5228_ VGND VPWR _0698_ _0605_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5159_ VPWR VGND VGND VPWR _0593_ _0629_ _3796_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_79_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_66_302 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_39_538 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_105_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_104_175 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_666 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_53_552 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4530_ VPWR VGND _4068_ round_key[69] new_block[69] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_104_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_4_159 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4461_ VGND VPWR _3999_ _3990_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6200_ _1437_ _1661_ _1288_ _1433_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7180_ VGND VPWR _2630_ _1198_ _2552_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6131_ VPWR VGND _1376_ _1592_ _1396_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_4392_ VGND VPWR _3930_ _3929_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_0_365 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6062_ VPWR VGND VGND VPWR _1524_ _1441_ _1375_ ZI_sky130_fd_sc_hd__nand2_2
X_5013_ VPWR VGND _0485_ _0301_ _0142_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_84_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_17_81 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_5_Right_5 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6964_ VPWR VGND _2417_ _2416_ _0447_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5915_ VPWR VGND VGND VPWR _3775_ _1377_ _1324_ _1329_ ZI_sky130_fd_sc_hd__nor3b_2
X_6895_ VGND VPWR VGND VPWR _2348_ _2344_ _2343_ _2346_ _2347_ ZI_sky130_fd_sc_hd__a211o_2
X_5846_ VPWR VGND VGND VPWR _1307_ _1308_ _1295_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_76_666 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5777_ VPWR VGND _1241_ new_block[110] round_key[110] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8496_ VGND VPWR VPWR VGND clk _0098_ reset_n new_block[55] ZI_sky130_fd_sc_hd__dfrtp_2
X_7516_ VPWR VGND VPWR VGND _2892_ _2948_ _2857_ _2880_ _4076_ _2949_ ZI_sky130_fd_sc_hd__a221o_2
X_4728_ VPWR VGND VGND VPWR _3965_ _0204_ _3804_ ZI_sky130_fd_sc_hd__nor2_2
X_4659_ VPWR VGND VGND VPWR _3962_ _3954_ _3999_ _3862_ _4196_ _4195_ ZI_sky130_fd_sc_hd__o221a_2
XFILLER_0_102_602 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7447_ VGND VPWR _2885_ _1997_ _2884_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_181 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_31_246 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7378_ VPWR VGND _2821_ _0986_ _0910_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_102_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6329_ VPWR VGND VGND VPWR _1479_ _1788_ _1609_ ZI_sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_103_Left_216 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_13_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_81_179 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_112_Left_225 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5700_ VGND VPWR VGND VPWR _0640_ _0652_ _1165_ _0783_ ZI_sky130_fd_sc_hd__a21oi_2
X_6680_ VPWR VGND _2113_ _2134_ _2133_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5631_ VPWR VGND VPWR VGND _1052_ _1096_ _1092_ _0945_ _1097_ ZI_sky130_fd_sc_hd__or4_2
X_5562_ VGND VPWR VGND VPWR _1029_ _0678_ _0929_ _0619_ ZI_sky130_fd_sc_hd__o21a_2
X_8350_ VGND VPWR VGND VPWR _3640_ new_block[26] _3705_ _3703_ _2483_ _0133_ ZI_sky130_fd_sc_hd__o32a_2
X_8281_ VGND VPWR _3643_ _2846_ _2849_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_533 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_53_371 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_53_393 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7301_ VPWR VGND VPWR VGND _2664_ _2128_ _2680_ _2229_ _2259_ _2748_ ZI_sky130_fd_sc_hd__a221o_2
X_4513_ VGND VPWR VPWR VGND _4049_ _4050_ _4048_ _4051_ ZI_sky130_fd_sc_hd__or3_2
X_7232_ VPWR VGND _2097_ _2681_ _2230_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5493_ VPWR VGND _0613_ _0961_ _0771_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_1_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4444_ VGND VPWR _3982_ _3849_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7163_ VGND VPWR VPWR VGND _2611_ _2612_ _2610_ _2613_ ZI_sky130_fd_sc_hd__or3_2
X_4375_ VGND VPWR _3913_ _3912_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7094_ VGND VPWR VPWR VGND _2515_ _2544_ _2504_ _2545_ ZI_sky130_fd_sc_hd__or3_2
X_6114_ VPWR VGND _1576_ _1575_ _1574_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6045_ VPWR VGND VPWR VGND _1414_ _1507_ _1313_ _1319_ ZI_sky130_fd_sc_hd__or3b_2
X_7996_ VPWR VGND _3385_ _0801_ _0799_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6947_ VGND VPWR VGND VPWR _2400_ _2157_ _2227_ _2189_ ZI_sky130_fd_sc_hd__o21a_2
X_6878_ VGND VPWR VPWR VGND _2331_ _2097_ _2168_ _2202_ _2231_ ZI_sky130_fd_sc_hd__o31a_2
XFILLER_0_63_113 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5829_ sword_ctr_reg\[1\] _1291_ sword_ctr_reg\[0\] new_block[17] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_91_444 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_8_284 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_44_360 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_106_259 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8479_ VGND VPWR VPWR VGND clk _0081_ reset_n new_block[38] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_12_290 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_40_59 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_54_168 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_105_281 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_50_396 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_4_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_65_23 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7850_ VGND VPWR _3253_ _2484_ _2559_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6801_ VGND VPWR _2255_ _2245_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4993_ VPWR VGND VPWR VGND _0457_ _0464_ _0460_ _0452_ _0465_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_105_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7781_ VGND VPWR _3190_ _1578_ _1680_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_430 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_260 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6732_ VGND VPWR _2186_ _2103_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_85_293 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6663_ VPWR VGND VGND VPWR _2078_ _2117_ _3850_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_5_221 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_45_146 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8402_ VPWR VGND VPWR VGND ready reset_n _0004_ clk ZI_sky130_fd_sc_hd__dfstp_2
XFILLER_0_61_617 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5614_ VGND VPWR VGND VPWR _1080_ _0757_ _0675_ _0717_ _0787_ _0923_ ZI_sky130_fd_sc_hd__a32o_2
X_6594_ VPWR VGND VPWR VGND _1281_ _1909_ _2048_ _1959_ _2047_ _2049_ ZI_sky130_fd_sc_hd__a221o_2
X_5545_ VGND VPWR VGND VPWR _0729_ _0661_ _0973_ _1012_ ZI_sky130_fd_sc_hd__a21o_2
X_8333_ VGND VPWR _3690_ _1830_ _3689_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8264_ VPWR VGND _3628_ block[50] round_key[50] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5476_ VGND VPWR VGND VPWR _0944_ _0589_ _0717_ _0601_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_76_3 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8195_ VGND VPWR VGND VPWR _3548_ new_block[11] _3565_ _3563_ _1054_ _0118_ ZI_sky130_fd_sc_hd__o32a_2
X_7215_ VGND VPWR VGND VPWR _2664_ _2135_ _2131_ _2119_ ZI_sky130_fd_sc_hd__o21a_2
X_4427_ VPWR VGND VPWR VGND _3891_ _3915_ _3932_ _3890_ _3965_ ZI_sky130_fd_sc_hd__or4_2
X_7146_ VGND VPWR VPWR VGND _2592_ _2595_ _2461_ _2596_ ZI_sky130_fd_sc_hd__or3_2
X_4358_ VGND VPWR _3896_ _3874_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7077_ VGND VPWR VGND VPWR _2528_ _2228_ _2368_ _2373_ ZI_sky130_fd_sc_hd__o21a_2
X_4289_ VGND VPWR VGND VPWR new_block[37] _3762_ _3825_ _3764_ _3827_ _3826_ ZI_sky130_fd_sc_hd__a221oi_2
X_6028_ VGND VPWR VPWR VGND _1333_ _1348_ _3796_ _1490_ ZI_sky130_fd_sc_hd__or3_2
X_7979_ VGND VPWR _3370_ _0153_ _3369_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_569 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_68_249 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_37_625 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_83_219 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_64_477 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_10_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_28_614 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_51_69 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_43_639 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_55_499 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5330_ VPWR VGND _0800_ round_key[46] new_block[46] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5261_ VPWR VGND VGND VPWR _0632_ _0731_ _0650_ ZI_sky130_fd_sc_hd__nor2_2
X_7000_ VPWR VGND VGND VPWR _2452_ _2174_ _2139_ ZI_sky130_fd_sc_hd__nand2_2
X_4212_ VPWR VGND VPWR VGND round[3] round[0] round[1] round[2] _3759_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_76_44 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5192_ VGND VPWR _0662_ _0661_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7902_ VGND VPWR VGND VPWR _3300_ _3299_ _3298_ _3296_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_92_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7833_ VPWR VGND _3238_ block[105] round_key[105] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_25_92 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7764_ VPWR VGND VGND VPWR _3174_ _3175_ _3170_ ZI_sky130_fd_sc_hd__nor2_2
X_6715_ VPWR VGND VGND VPWR _2147_ _2169_ _2110_ ZI_sky130_fd_sc_hd__nor2_2
X_4976_ VGND VPWR VGND VPWR _4104_ new_block[101] _0448_ _0445_ _0429_ _0016_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_46_477 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7695_ VGND VPWR _3112_ _0232_ _0311_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_105 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6646_ VGND VPWR VGND VPWR _2064_ _3914_ _2100_ _2063_ ZI_sky130_fd_sc_hd__nand3_2
X_6577_ VGND VPWR VGND VPWR _1614_ _1534_ _1480_ _2032_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_104_527 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5528_ VPWR VGND _0996_ _0811_ _0806_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8316_ VGND VPWR VPWR VGND _3673_ _3669_ _3675_ _0366_ _3674_ ZI_sky130_fd_sc_hd__o211a_2
X_8247_ VGND VPWR VGND VPWR _3548_ new_block[16] _3612_ _3610_ _1562_ _0123_ ZI_sky130_fd_sc_hd__o32a_2
X_5459_ VGND VPWR VPWR VGND _0596_ _0926_ _0925_ _0927_ ZI_sky130_fd_sc_hd__mux2_2
X_8178_ VGND VPWR _3550_ _0381_ _3549_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7129_ VPWR VGND _2345_ _2579_ _2173_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_37_466 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_25_639 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_37_488 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_92_583 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_1_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4830_ VPWR VGND _0305_ round_key[66] new_block[66] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4761_ VGND VPWR _0237_ _0233_ _0236_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_349 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6500_ VGND VPWR VGND VPWR _1956_ _1954_ _1957_ _1001_ ZI_sky130_fd_sc_hd__a21oi_2
X_7480_ VPWR VGND _2915_ _1751_ _1683_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4692_ VGND VPWR _0169_ _0168_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_102_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6431_ VPWR VGND _1889_ _1888_ _1682_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_11_94 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_102_85 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6362_ VGND VPWR _1821_ _1568_ _1820_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5313_ VPWR VGND VGND VPWR _0783_ _0583_ _0609_ ZI_sky130_fd_sc_hd__nand2_2
X_8101_ VPWR VGND VPWR VGND _3459_ _3367_ _3480_ _3468_ _1751_ _3481_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_3_599 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6293_ VGND VPWR _1753_ _1566_ _1688_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8032_ VPWR VGND _3418_ _1132_ _1131_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5244_ VPWR VGND _0683_ _0714_ _0713_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5175_ VGND VPWR _0645_ _0644_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7816_ VGND VPWR _3222_ _2558_ _3221_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_444 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4959_ VPWR VGND _0432_ _0431_ _0367_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7747_ VPWR VGND VPWR VGND _3150_ _3159_ _3158_ _3139_ _0908_ _3160_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_19_477 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7678_ VPWR VGND _3096_ _0431_ _0370_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6629_ VGND VPWR VGND VPWR _2083_ _3822_ _2079_ _2080_ _2081_ _2082_ ZI_sky130_fd_sc_hd__a41o_2
XFILLER_0_14_160 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_97_642 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_96_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_69_377 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_65_561 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_52_211 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_57_46 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6980_ VGND VPWR VGND VPWR _2432_ _2162_ _2182_ _2252_ _2118_ ZI_sky130_fd_sc_hd__and4_2
X_5931_ VPWR VGND VGND VPWR _1393_ _3914_ _1392_ ZI_sky130_fd_sc_hd__nand2_2
X_5862_ VGND VPWR VGND VPWR _3797_ _1320_ _1321_ _1322_ _1324_ _1323_ ZI_sky130_fd_sc_hd__o41ai_2
XFILLER_0_87_196 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_8_614 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4813_ VPWR VGND VGND VPWR _0288_ _0287_ _0286_ _4164_ _4025_ _3955_ ZI_sky130_fd_sc_hd__o2111a_2
X_5793_ VGND VPWR VGND VPWR _1256_ _0859_ _0787_ _0628_ _0975_ _0923_ ZI_sky130_fd_sc_hd__a32o_2
X_7601_ VGND VPWR _3026_ _0319_ _2687_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4744_ VGND VPWR VPWR VGND _3982_ _3862_ _0220_ _0219_ _0217_ ZI_sky130_fd_sc_hd__o211a_2
X_7532_ VGND VPWR _2963_ _2004_ _2962_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_22_71 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4675_ VPWR VGND _0152_ round_key[81] new_block[81] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_98_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7463_ VGND VPWR VPWR VGND _2898_ _2897_ _2900_ _2855_ _2899_ ZI_sky130_fd_sc_hd__o211a_2
X_7394_ VGND VPWR _2836_ _1229_ _2835_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6414_ VGND VPWR VGND VPWR _1653_ _1538_ _1399_ _1436_ _1344_ _1872_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_43_299 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6345_ _1515_ _1804_ _1334_ _1409_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6276_ _1734_ _1736_ _1733_ _1735_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8015_ VPWR VGND VPWR VGND _3309_ _3367_ _3402_ _3328_ _0988_ _3403_ ZI_sky130_fd_sc_hd__a221o_2
X_5227_ VGND VPWR VPWR VGND _0695_ _0696_ _0658_ _0697_ ZI_sky130_fd_sc_hd__or3_2
X_5158_ VGND VPWR _0628_ _0627_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_98_417 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5089_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] _0559_ new_block[78] ZI_sky130_fd_sc_hd__and2b_2
XFILLER_0_79_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_94_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_78_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_78_174 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_47_561 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_22_428 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_104_187 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_27_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_89_428 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_43_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_72_317 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_5_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_25_233 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_25_244 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_7_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4460_ VGND VPWR _3998_ _3971_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4391_ VGND VPWR VPWR VGND _3809_ _3814_ _3850_ _3929_ ZI_sky130_fd_sc_hd__or3_2
X_6130_ VGND VPWR VGND VPWR _1591_ _1511_ _1337_ _1589_ _1590_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_0_355 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_0_377 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6061_ VGND VPWR _1523_ _1408_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5012_ VGND VPWR _0484_ _0479_ _0483_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6963_ VGND VPWR _2416_ _0164_ _0489_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5914_ _1335_ _1376_ _1334_ _1375_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6894_ VGND VPWR VGND VPWR _2347_ _2174_ _2282_ _2115_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_76_645 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_8_411 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5845_ VGND VPWR _1307_ _1306_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_75_122 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_29_561 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5776_ VPWR VGND _1240_ block[46] round_key[46] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_44_542 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8495_ VGND VPWR VPWR VGND clk _0097_ reset_n new_block[54] ZI_sky130_fd_sc_hd__dfrtp_2
X_7515_ VPWR VGND _2948_ block[13] round_key[13] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4727_ VGND VPWR VGND VPWR _4134_ _3817_ _3982_ _3895_ _0203_ ZI_sky130_fd_sc_hd__a2bb2o_2
X_4658_ VGND VPWR VGND VPWR _3872_ _3918_ _4023_ _3990_ _4195_ ZI_sky130_fd_sc_hd__o22a_2
X_7446_ VPWR VGND _2884_ _1577_ _1574_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_3_160 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_101_113 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_102_614 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_101_146 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7377_ VGND VPWR VGND VPWR _2800_ new_block[66] _2820_ _2818_ _0229_ _0045_ ZI_sky130_fd_sc_hd__o32a_2
X_4589_ VGND VPWR VGND VPWR _4125_ _3816_ _4126_ _3990_ ZI_sky130_fd_sc_hd__a21oi_2
X_6328_ VPWR VGND VPWR VGND _1700_ _1786_ _1785_ _1536_ _1787_ ZI_sky130_fd_sc_hd__or4_2
X_6259_ VPWR VGND VPWR VGND _1588_ _1719_ _1368_ _1462_ ZI_sky130_fd_sc_hd__or3b_2
XPHY_EDGE_ROW_11_Right_11 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_66_133 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_66_177 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_35_575 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_50_578 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_50_589 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_20_Right_20 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_85_475 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_73_637 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_70_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_57_188 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5630_ VGND VPWR VGND VPWR _1093_ _0532_ _0949_ _1094_ _1096_ _1095_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_26_564 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_41_501 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5561_ VPWR VGND VPWR VGND _1027_ _0639_ _1025_ _0722_ _1024_ _1028_ ZI_sky130_fd_sc_hd__a221o_2
X_8280_ VGND VPWR _3642_ _0914_ _3641_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_225 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_53_383 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7300_ VGND VPWR VGND VPWR _2229_ _2338_ _2437_ _2501_ _2747_ _2516_ ZI_sky130_fd_sc_hd__a2111o_2
X_5492_ VPWR VGND VPWR VGND _0959_ _0847_ _0674_ _0653_ _0960_ ZI_sky130_fd_sc_hd__a22o_2
X_4512_ VGND VPWR VGND VPWR _4036_ _3971_ _4050_ _3859_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_41_545 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7231_ VPWR VGND _2190_ _2680_ _2368_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_110_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_1_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_110_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4443_ VPWR VGND VGND VPWR _3887_ _3981_ _3895_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_0_141 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7162_ VPWR VGND VPWR VGND _2173_ _2368_ _2120_ _2135_ _2612_ ZI_sky130_fd_sc_hd__a22o_2
X_4374_ VGND VPWR VGND VPWR _3912_ _3846_ _3837_ _3885_ ZI_sky130_fd_sc_hd__and3b_2
X_7093_ VPWR VGND VPWR VGND _2537_ _2543_ _2539_ _2530_ _2544_ ZI_sky130_fd_sc_hd__or4_2
X_6113_ VPWR VGND _1575_ round_key[24] new_block[24] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6044_ _1331_ _1506_ _1288_ _1437_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_21_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7995_ VGND VPWR VGND VPWR _3331_ new_block[56] _3384_ _3382_ _2307_ _0099_ ZI_sky130_fd_sc_hd__o32a_2
X_6946_ VPWR VGND VPWR VGND _2157_ _2215_ _2195_ _2170_ _2399_ ZI_sky130_fd_sc_hd__a22o_2
X_6877_ VGND VPWR _2330_ _2264_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5828_ VGND VPWR VGND VPWR _1290_ new_block[49] sword_ctr_reg\[1\] sword_ctr_reg\[0\]
+ ZI_sky130_fd_sc_hd__and3b_2
X_5759_ VGND VPWR VGND VPWR _0645_ _0675_ _0978_ _0877_ _1223_ _0867_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_63_169 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_32_567 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8478_ VGND VPWR VPWR VGND clk _0080_ reset_n new_block[37] ZI_sky130_fd_sc_hd__dfrtp_2
X_7429_ VGND VPWR _2869_ _2865_ _2868_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_86_239 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_94_261 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_67_486 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_2_417 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_65_57 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6800_ VPWR VGND VPWR VGND _2253_ _2131_ _2213_ _2148_ _2245_ _2254_ ZI_sky130_fd_sc_hd__a221o_2
X_4992_ VPWR VGND VPWR VGND _0463_ _0464_ _0461_ _0462_ ZI_sky130_fd_sc_hd__or3b_2
X_7780_ VGND VPWR _3189_ _1574_ _1885_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6731_ VGND VPWR VGND VPWR _2185_ _2184_ _2149_ _2144_ ZI_sky130_fd_sc_hd__o21a_2
X_6662_ VPWR VGND _2112_ _2116_ _2115_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5613_ _0648_ _1079_ _0704_ _0851_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_45_169 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8401_ VGND VPWR VPWR VGND clk _0001_ reset_n dec_ctrl_reg\[3\] ZI_sky130_fd_sc_hd__dfrtp_2
X_6593_ VPWR VGND _2048_ new_block[119] round_key[119] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8332_ VGND VPWR _3689_ _1576_ _3688_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5544_ VPWR VGND VPWR VGND _1010_ _0929_ _0771_ _0602_ _0712_ _1011_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_103_208 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8263_ VGND VPWR VGND VPWR _3627_ _3626_ _3625_ _3621_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_14_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5475_ VPWR VGND VPWR VGND _0588_ _0751_ _0746_ _0739_ _0943_ ZI_sky130_fd_sc_hd__a22o_2
X_4426_ VPWR VGND VGND VPWR _3964_ _3958_ _3963_ ZI_sky130_fd_sc_hd__nand2_2
X_8194_ VPWR VGND VPWR VGND _3459_ _3490_ _3564_ _3468_ _1816_ _3565_ ZI_sky130_fd_sc_hd__a221o_2
X_7214_ VGND VPWR VGND VPWR _2663_ _2658_ _2343_ _2659_ _2662_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_111_263 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_69_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7145_ VGND VPWR VPWR VGND _2519_ _2594_ _2593_ _2595_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_39_80 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4357_ VPWR VGND VGND VPWR _3895_ _3894_ _3795_ ZI_sky130_fd_sc_hd__nand2_2
X_7076_ VGND VPWR VGND VPWR _2526_ _2525_ _2173_ _2139_ _2527_ ZI_sky130_fd_sc_hd__a31o_2
X_4288_ sword_ctr_reg\[1\] _3826_ sword_ctr_reg\[0\] new_block[5] VPWR VGND VPWR VGND
+ ZI_sky130_fd_sc_hd__and3_2
X_6027_ _1319_ _1489_ _1313_ _1414_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7978_ VGND VPWR _3369_ _0383_ _0514_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6929_ VPWR VGND VPWR VGND _2382_ _3776_ _2094_ ZI_sky130_fd_sc_hd__or2_2
XFILLER_0_9_561 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_37_637 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_20_559 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_102_263 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_121 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_19_39 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_95_570 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_27_169 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_2_247 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5260_ VGND VPWR VGND VPWR _0730_ _0727_ _0726_ _0589_ _0729_ _0655_ ZI_sky130_fd_sc_hd__a32o_2
X_4211_ VPWR VGND VGND VPWR _0001_ _3758_ _0000_ ZI_sky130_fd_sc_hd__nor2_2
X_5191_ VGND VPWR _0661_ _0656_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_76_56 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7901_ VGND VPWR VGND VPWR _3298_ _3296_ _3299_ _3028_ ZI_sky130_fd_sc_hd__a21oi_2
X_7832_ VGND VPWR _3237_ _2702_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7763_ VGND VPWR _3174_ _3172_ _3173_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4975_ VPWR VGND VPWR VGND _4101_ _0169_ _0447_ _0162_ _0446_ _0448_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_18_103 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6714_ VGND VPWR _2168_ _2167_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_73_220 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_18_158 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_46_445 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7694_ VGND VPWR _3111_ _0142_ _0301_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_46_489 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6645_ VPWR VGND VGND VPWR _2099_ _3914_ _2098_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_61_437 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6576_ VGND VPWR VGND VPWR _1506_ _1395_ _1368_ _1434_ _2031_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_42_640 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5527_ VGND VPWR _0995_ _0992_ _0994_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8315_ VPWR VGND VGND VPWR _3674_ _3669_ _3673_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_41_150 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8246_ VPWR VGND VPWR VGND _3575_ _3603_ _3611_ _3583_ _1676_ _3612_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_112_561 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5458_ VPWR VGND VGND VPWR _0926_ _0580_ _0571_ ZI_sky130_fd_sc_hd__nand2_2
X_4409_ _3945_ _3947_ _3795_ _3946_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8177_ VPWR VGND _3549_ _0155_ _4077_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5389_ VGND VPWR VGND VPWR _0850_ _0639_ _0853_ _0855_ _0858_ _0857_ ZI_sky130_fd_sc_hd__a2111o_2
X_7128_ VGND VPWR VGND VPWR _2578_ _2378_ _2166_ _2268_ _2266_ ZI_sky130_fd_sc_hd__a211o_2
X_7059_ VPWR VGND VPWR VGND _2327_ _2194_ _2107_ _2302_ _2510_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_37_445 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_103_561 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_87_301 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4760_ VGND VPWR _0236_ _0234_ _0235_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_112_Right_112 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4691_ VGND VPWR _0168_ _0167_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_11_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_102_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6430_ VGND VPWR _1888_ _1571_ _1759_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6361_ VPWR VGND _1820_ round_key[18] new_block[18] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_30_109 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8100_ VPWR VGND _3480_ block[98] round_key[98] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5312_ VPWR VGND VPWR VGND _0781_ _0532_ _0779_ _0596_ _0778_ _0782_ ZI_sky130_fd_sc_hd__a221o_2
X_6292_ VGND VPWR _1752_ _1563_ _1751_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8031_ VGND VPWR _3417_ _1130_ _3416_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5243_ VPWR VGND _0581_ _0713_ _0586_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5174_ _0642_ _0644_ _0581_ _0643_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_58_Right_58 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7815_ VPWR VGND _3221_ _2411_ _2316_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_109_609 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_59_581 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4958_ VPWR VGND _0431_ round_key[68] new_block[68] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7746_ VGND VPWR _3159_ _0161_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7677_ VPWR VGND _3095_ _0436_ _0155_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4889_ VGND VPWR _0363_ new_block[100] round_key[100] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_89_Left_202 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6628_ VPWR VGND VGND VPWR sword_ctr_reg\[0\] sword_ctr_reg\[1\] new_block[120] _2082_
+ ZI_sky130_fd_sc_hd__nor3_2
XPHY_EDGE_ROW_67_Right_67 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6559_ VGND VPWR VGND VPWR _2014_ _1478_ _1390_ _1988_ _2013_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_14_172 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_30_610 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_42_492 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_100_520 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_100_542 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8229_ VGND VPWR _3596_ _0435_ _3123_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_98_Left_211 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Right_76 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_97_654 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_65_573 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_85_Right_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_110_328 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Right_94 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5930_ VGND VPWR VPWR VGND _1303_ _1302_ _1301_ _4097_ _1304_ _1392_ ZI_sky130_fd_sc_hd__a41oi_2
XFILLER_0_73_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5861_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[117] sword_ctr_reg\[0\] _1323_
+ ZI_sky130_fd_sc_hd__or3_2
X_7600_ VGND VPWR _3025_ _3021_ _3024_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_103 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_8_626 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4812_ VGND VPWR VGND VPWR _4016_ _3918_ _3933_ _0287_ ZI_sky130_fd_sc_hd__a21o_2
X_5792_ VGND VPWR VPWR VGND _1252_ _1254_ _1250_ _1255_ ZI_sky130_fd_sc_hd__or3_2
X_4743_ VPWR VGND VGND VPWR _0219_ _4030_ _0218_ ZI_sky130_fd_sc_hd__nand2_2
X_7531_ VPWR VGND _2962_ _1997_ _1898_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_7_169 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7462_ VPWR VGND VGND VPWR _2899_ _2897_ _2898_ ZI_sky130_fd_sc_hd__nand2_2
X_6413_ VGND VPWR VPWR VGND _1405_ _1436_ _1344_ _1871_ ZI_sky130_fd_sc_hd__or3_2
X_4674_ VGND VPWR _0151_ _0148_ _0150_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7393_ VGND VPWR _2835_ _0805_ _1069_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6344_ VPWR VGND VPWR VGND _1802_ _1376_ _1639_ _1511_ _1604_ _1803_ ZI_sky130_fd_sc_hd__a221o_2
X_6275_ VGND VPWR VGND VPWR _1475_ _1445_ _1384_ _1735_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_11_197 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8014_ VPWR VGND _3402_ block[58] round_key[58] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5226_ _0577_ _0696_ _0630_ _0579_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_51_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5157_ VPWR VGND _0605_ _0627_ _0626_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5088_ VGND VPWR VGND VPWR _0558_ new_block[46] sword_ctr_reg\[1\] sword_ctr_reg\[0\]
+ ZI_sky130_fd_sc_hd__and3b_2
XFILLER_0_79_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_94_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_109_406 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_47_573 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7729_ VGND VPWR _3143_ _1825_ _3142_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_576 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_15_470 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_34_278 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_62_598 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_27_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_57_304 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_57_337 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_5_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_40_204 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4390_ VGND VPWR VPWR VGND _3922_ _3927_ _3919_ _3928_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_0_389 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6060_ VGND VPWR _1522_ _1379_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5011_ VGND VPWR _0483_ _0481_ _0482_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_108_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6962_ VPWR VGND _2415_ _2414_ _2410_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_76_602 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5913_ VGND VPWR VGND VPWR _1294_ _1347_ _3796_ _1375_ ZI_sky130_fd_sc_hd__a21o_2
X_6893_ _2345_ _2346_ _2118_ _2199_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_75_101 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5844_ VGND VPWR VPWR VGND _1300_ _1305_ _3787_ _1306_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_29_573 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_33_93 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5775_ VGND VPWR VPWR VGND _1237_ _1231_ _1239_ _0444_ _1238_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_99_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7514_ VGND VPWR VGND VPWR _2947_ _2946_ _2945_ _2943_ ZI_sky130_fd_sc_hd__o21a_2
X_8494_ VGND VPWR VPWR VGND clk _0096_ reset_n new_block[53] ZI_sky130_fd_sc_hd__dfrtp_2
X_4726_ VPWR VGND VPWR VGND _4159_ _0201_ _0199_ _4024_ _0202_ ZI_sky130_fd_sc_hd__or4_2
X_4657_ VPWR VGND VPWR VGND _4191_ _4193_ _4194_ _4187_ _4190_ ZI_sky130_fd_sc_hd__or4b_2
X_7445_ VPWR VGND _2883_ _1680_ _1575_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_102_626 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7376_ VPWR VGND VPWR VGND _2797_ _2786_ _2819_ _2703_ _0305_ _2820_ ZI_sky130_fd_sc_hd__a221o_2
X_6327_ VPWR VGND VPWR VGND _1491_ _1493_ _1437_ _1426_ _1786_ ZI_sky130_fd_sc_hd__a22o_2
X_4588_ VPWR VGND VGND VPWR _4125_ _3878_ _3868_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_101_169 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6258_ VGND VPWR VGND VPWR _1717_ _1521_ _1718_ _1716_ ZI_sky130_fd_sc_hd__a21bo_2
X_6189_ VGND VPWR _1427_ _1421_ _1650_ _1604_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
X_5209_ VGND VPWR VGND VPWR _0679_ _0669_ _0675_ _0651_ _0678_ _0674_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_39_337 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_109_225 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_47_381 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_82_638 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_81_126 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_26_Left_139 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_54_15 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_54_48 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_54_59 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_35_Left_148 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_97_281 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_70_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_57_156 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_73_649 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5560_ VPWR VGND VPWR VGND _1026_ _0717_ _0702_ _0706_ _0751_ _1027_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_26_576 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5491_ VPWR VGND VPWR VGND _0959_ _3777_ _0537_ ZI_sky130_fd_sc_hd__or2_2
X_4511_ VPWR VGND VPWR VGND _3869_ _3924_ _3845_ _3923_ _4049_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_1_610 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4442_ VPWR VGND VPWR VGND _3972_ _3979_ _3977_ _3968_ _3980_ ZI_sky130_fd_sc_hd__or4_2
X_7230_ VPWR VGND VPWR VGND _2284_ _2249_ _2679_ _2340_ _2295_ ZI_sky130_fd_sc_hd__or4b_2
XFILLER_0_110_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Left_157 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_111_445 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_0_153 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_1_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_21_281 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_110_97 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7161_ VGND VPWR VGND VPWR _2611_ _2231_ _2297_ _2120_ _2259_ _2207_ ZI_sky130_fd_sc_hd__a32o_2
X_4373_ VPWR VGND VGND VPWR _3910_ _3911_ _3877_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_0_197 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6112_ VPWR VGND _1574_ round_key[29] new_block[29] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7092_ VGND VPWR VGND VPWR _2299_ _2203_ _2294_ _2541_ _2543_ _2542_ ZI_sky130_fd_sc_hd__a2111o_2
X_6043_ VPWR VGND VPWR VGND _1500_ _1504_ _1502_ _1497_ _1505_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_95_99 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7994_ VPWR VGND VPWR VGND _3309_ _3367_ _3383_ _3328_ _0806_ _3384_ ZI_sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_53_Left_166 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_49_602 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6945_ VGND VPWR VGND VPWR _2398_ _2278_ _2182_ _2173_ _2239_ _2397_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_44_81 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_49_635 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6876_ VPWR VGND VPWR VGND _2325_ _2225_ _2326_ _2328_ _2329_ ZI_sky130_fd_sc_hd__or4bb_2
XFILLER_0_8_253 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5827_ VGND VPWR _1289_ _1288_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_76_498 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_8_297 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5758_ VGND VPWR VGND VPWR _0741_ _0677_ _1221_ _0873_ _1222_ _0970_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_32_513 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4709_ _3838_ _0185_ _3831_ _3901_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8477_ VGND VPWR VPWR VGND clk _0079_ reset_n new_block[36] ZI_sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_62_Left_175 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7428_ VGND VPWR _2868_ _2866_ _2867_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_181 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5689_ _0689_ _1154_ _0674_ _0787_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_32_579 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7359_ VGND VPWR _2804_ _2788_ _2803_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_71_Left_184 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_24_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_86_218 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_39_178 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_67_498 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_80_Left_193 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_23_524 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_112_209 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_105_294 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4991_ VGND VPWR VGND VPWR _3976_ _4125_ _4116_ _4141_ _0463_ ZI_sky130_fd_sc_hd__o22a_2
X_6730_ VGND VPWR _2184_ _2183_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_81_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_273 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6661_ VGND VPWR _2115_ _2114_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6592_ VPWR VGND _2047_ block[23] round_key[23] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5612_ VGND VPWR VGND VPWR _1009_ new_block[107] _1078_ _1056_ _1054_ _0022_ ZI_sky130_fd_sc_hd__o32a_2
X_8400_ VGND VPWR VPWR VGND clk _0000_ reset_n dec_ctrl_reg\[2\] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_245 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5543_ VPWR VGND VPWR VGND _0701_ _0692_ _0589_ _0658_ _1010_ ZI_sky130_fd_sc_hd__a22o_2
X_8331_ VGND VPWR _3688_ _1578_ _3687_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_332 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_53_181 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8262_ VGND VPWR VGND VPWR _3625_ _3621_ _3626_ _4085_ ZI_sky130_fd_sc_hd__a21oi_2
X_5474_ _0618_ _0942_ _0687_ _0677_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_4425_ VGND VPWR VGND VPWR _3930_ _3906_ _3962_ _3959_ _3932_ _3963_ ZI_sky130_fd_sc_hd__o32a_2
X_7213_ VPWR VGND VPWR VGND _2224_ _2661_ _2660_ _2217_ _2662_ ZI_sky130_fd_sc_hd__or4_2
X_8193_ VPWR VGND _3564_ block[75] round_key[75] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4356_ VGND VPWR VGND VPWR _3814_ _3809_ _3776_ _3894_ ZI_sky130_fd_sc_hd__a21o_2
X_7144_ VGND VPWR VGND VPWR _2594_ _2222_ _2236_ _2112_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_39_92 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7075_ VPWR VGND VGND VPWR _2526_ _2175_ _2163_ _2139_ _2138_ _2162_ ZI_sky130_fd_sc_hd__o2111a_2
X_4287_ VPWR VGND VGND VPWR new_block[69] sword_ctr_reg\[0\] _3825_ ZI_sky130_fd_sc_hd__or2b_2
X_6026_ VGND VPWR VGND VPWR _1473_ _1466_ _1488_ _1487_ ZI_sky130_fd_sc_hd__a21oi_2
X_7977_ VGND VPWR VGND VPWR _3331_ new_block[54] _3368_ _3365_ _1996_ _0097_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_49_465 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6928_ VPWR VGND VPWR VGND _2102_ _2131_ _2123_ _2173_ _2381_ ZI_sky130_fd_sc_hd__a22o_2
X_6859_ VGND VPWR _2313_ _2309_ _2312_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_37_649 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_32_332 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8529_ VGND VPWR VPWR VGND clk _0131_ reset_n new_block[24] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_72_490 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_32_365 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_102_253 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_3_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_102_275 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_87_505 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_109_Left_222 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_82_221 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_67_262 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_55_468 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_35_192 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_51_663 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4210_ VGND VPWR _0001_ _3757_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5190_ VGND VPWR VGND VPWR _0660_ _0651_ _0648_ _0653_ _0659_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_76_68 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7900_ VGND VPWR _3298_ _3084_ _3297_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7831_ VGND VPWR VGND VPWR _3236_ _3235_ _3234_ _3230_ ZI_sky130_fd_sc_hd__o21a_2
X_7762_ VPWR VGND _3173_ _1830_ _1763_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4974_ VPWR VGND _0447_ new_block[101] round_key[101] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7693_ VGND VPWR _3110_ _3107_ _3109_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6713_ VPWR VGND _2129_ _2167_ _2166_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_46_457 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6644_ VGND VPWR VGND VPWR _0538_ _2065_ _2066_ _2067_ _2068_ _2098_ ZI_sky130_fd_sc_hd__o41a_2
X_6575_ VPWR VGND VPWR VGND _1698_ _1515_ _1546_ _1527_ _1434_ _2030_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_14_321 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_26_192 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_33_129 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_81_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5526_ VPWR VGND _0994_ _0993_ _0912_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_14_365 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8314_ VGND VPWR _3673_ _3671_ _3672_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8245_ VPWR VGND _3611_ block[48] round_key[48] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5457_ VPWR VGND VGND VPWR _0925_ _0846_ _0654_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_112_573 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4408_ VPWR VGND VGND VPWR _3890_ _3838_ _3885_ _3946_ ZI_sky130_fd_sc_hd__nor3_2
X_8176_ VGND VPWR VGND VPWR _3548_ new_block[9] _3547_ _3545_ _0899_ _0116_ ZI_sky130_fd_sc_hd__o32a_2
X_5388_ VGND VPWR VGND VPWR _0857_ _0780_ _0723_ _0652_ _0856_ _0584_ ZI_sky130_fd_sc_hd__o221ai_2
X_4339_ VGND VPWR _3877_ _3876_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7127_ VGND VPWR VGND VPWR _2577_ _2378_ _2339_ _2575_ _2576_ ZI_sky130_fd_sc_hd__a211o_2
X_7058_ VGND VPWR VPWR VGND _2507_ _2508_ _2234_ _2509_ ZI_sky130_fd_sc_hd__or3_2
X_6009_ _1335_ _1471_ _1334_ _1367_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_69_505 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_64_210 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_37_457 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_24_129 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_107_356 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_32_151 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_103_573 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_46_16 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_16_608 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4690_ _0166_ _0167_ _3749_ _3767_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_102_65 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6360_ VPWR VGND _1819_ round_key[27] new_block[27] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_3_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5311_ VGND VPWR VGND VPWR _0780_ _0774_ _0781_ _0640_ ZI_sky130_fd_sc_hd__a21oi_2
X_8030_ VGND VPWR _3416_ _1136_ _3415_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6291_ VPWR VGND _1751_ round_key[2] new_block[2] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5242_ VGND VPWR _0712_ _0711_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_87_78 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5173_ VGND VPWR VPWR VGND _0603_ _0604_ _3832_ _0643_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_78_324 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_93_305 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7814_ VGND VPWR VGND VPWR _3153_ new_block[39] _3220_ _3217_ _0513_ _0082_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_59_593 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_46_210 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7745_ VPWR VGND _3158_ block[1] round_key[1] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4957_ VGND VPWR _0430_ _4067_ _0305_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4888_ VGND VPWR VPWR VGND _0362_ _4123_ _0334_ _0361_ _3756_ ZI_sky130_fd_sc_hd__o31a_2
X_7676_ VGND VPWR VGND VPWR _2997_ new_block[91] _3094_ _3092_ _2545_ _0070_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_74_596 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6627_ VGND VPWR VGND VPWR sword_ctr_reg\[1\] sword_ctr_reg\[0\] new_block[88] _2081_
+ ZI_sky130_fd_sc_hd__nand3b_2
X_6558_ VGND VPWR VGND VPWR _2013_ _1639_ _1443_ _1727_ _1632_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_15_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5509_ VPWR VGND VPWR VGND _0976_ _0616_ _0710_ _0975_ _0702_ _0977_ ZI_sky130_fd_sc_hd__a221o_2
X_6489_ VGND VPWR _1946_ _1570_ _1945_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8228_ VGND VPWR VGND VPWR _3548_ new_block[14] _3595_ _3593_ _1227_ _0121_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_100_554 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8159_ VGND VPWR VGND VPWR _3462_ new_block[7] _3533_ _3529_ _0513_ _0114_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_97_611 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_97_666 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_32_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_65_541 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_65_585 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_80_533 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_60_290 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_103_370 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_73_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5860_ VGND VPWR VGND VPWR _1322_ sword_ctr_reg\[0\] new_block[85] sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__and3b_2
XFILLER_0_87_143 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4811_ VGND VPWR VGND VPWR _3916_ _3865_ _3854_ _0286_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_8_638 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5791_ VGND VPWR VGND VPWR _1254_ _0771_ _0859_ _1253_ _0636_ ZI_sky130_fd_sc_hd__a211o_2
X_4742_ VPWR VGND VGND VPWR _3910_ _0218_ _3930_ ZI_sky130_fd_sc_hd__nor2_2
X_7530_ VGND VPWR VGND VPWR _2894_ new_block[78] _2961_ _2958_ _1227_ _0057_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_71_500 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_56_585 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4673_ VGND VPWR _0150_ _4072_ _0149_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7461_ VGND VPWR _2898_ _1831_ _2887_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6412_ VGND VPWR _1390_ _1869_ _1870_ _1704_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
X_7392_ VPWR VGND _2834_ _2833_ _0909_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6343_ VPWR VGND VPWR VGND _1456_ _1419_ _1361_ _1408_ _1802_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_98_99 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6274_ VGND VPWR VGND VPWR _1412_ _1507_ _1371_ _1447_ _1734_ ZI_sky130_fd_sc_hd__o22a_2
X_8013_ VGND VPWR VGND VPWR _3401_ _3400_ _3399_ _3396_ ZI_sky130_fd_sc_hd__o21a_2
X_5225_ VGND VPWR _0695_ _0692_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_44_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5156_ VGND VPWR _0626_ _0587_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_47_81 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5087_ VPWR VGND VGND VPWR _0551_ _0555_ _0556_ _3914_ _0557_ ZI_sky130_fd_sc_hd__and4b_2
XFILLER_0_94_625 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_93_113 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_93_102 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_78_165 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5989_ VPWR VGND VPWR VGND _1387_ _1450_ _1411_ _1374_ _1451_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_93_135 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7728_ VPWR VGND _3142_ _1677_ _1570_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_47_585 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7659_ VGND VPWR _3079_ _3075_ _3078_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_181 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_108_473 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_80_341 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_40_216 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5010_ VPWR VGND _0482_ _0312_ _0153_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_108_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_17_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6961_ VGND VPWR _2414_ _2411_ _2413_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5912_ VGND VPWR VPWR VGND _1356_ _1373_ _1342_ _1374_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_48_305 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6892_ VGND VPWR _2345_ _2072_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5843_ VGND VPWR VGND VPWR _1305_ _3822_ _1301_ _1302_ _1303_ _1304_ ZI_sky130_fd_sc_hd__a41o_2
XFILLER_0_91_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5774_ VPWR VGND VGND VPWR _1238_ _1231_ _1237_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_29_585 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7513_ VGND VPWR VGND VPWR _2945_ _2943_ _2946_ _2642_ ZI_sky130_fd_sc_hd__a21oi_2
X_8493_ VGND VPWR VPWR VGND clk _0095_ reset_n new_block[52] ZI_sky130_fd_sc_hd__dfrtp_2
X_4725_ VGND VPWR VGND VPWR _0200_ _3898_ _3945_ _4010_ _0201_ ZI_sky130_fd_sc_hd__a31o_2
X_4656_ VGND VPWR VGND VPWR _4125_ _4036_ _3941_ _4192_ _4193_ ZI_sky130_fd_sc_hd__o22a_2
X_7444_ VGND VPWR VGND VPWR _2800_ new_block[71] _2882_ _2879_ _0513_ _0050_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_101_104 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7375_ VPWR VGND _2819_ block[34] round_key[34] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4587_ VGND VPWR VGND VPWR _3974_ _3859_ _4124_ _4036_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_3_195 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6326_ VPWR VGND VPWR VGND _1443_ _1419_ _1379_ _1408_ _1785_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_102_638 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6257_ VGND VPWR VGND VPWR _1524_ _1399_ _1473_ _1547_ _1424_ _1717_ ZI_sky130_fd_sc_hd__o32a_2
X_6188_ VGND VPWR _1511_ _1346_ _1649_ _1421_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
X_5208_ VGND VPWR _0678_ _0677_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5139_ VGND VPWR _0609_ _0608_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_39_327 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_109_237 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_35_533 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_35_588 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_105_432 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_70_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_57_135 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_73_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_499 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_53_352 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4510_ VPWR VGND _4046_ _4048_ _4047_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5490_ VPWR VGND VGND VPWR _0837_ _0958_ _0783_ ZI_sky130_fd_sc_hd__nor2_2
X_4441_ VGND VPWR VGND VPWR _3978_ _3954_ _3979_ _3962_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_102_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_110_65 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7160_ VGND VPWR VGND VPWR _2255_ _2202_ _2609_ _2610_ ZI_sky130_fd_sc_hd__a21o_2
X_6111_ VGND VPWR _1573_ _1567_ _1572_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4372_ VGND VPWR VGND VPWR _3802_ _3793_ _3910_ _3880_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_165 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7091_ VGND VPWR VGND VPWR _2542_ _2202_ _2231_ _2338_ ZI_sky130_fd_sc_hd__o21a_2
X_6042_ VGND VPWR VGND VPWR _1504_ _1397_ _1444_ _1390_ _1503_ _1336_ ZI_sky130_fd_sc_hd__a32o_2
XPHY_EDGE_ROW_107_Right_107 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7993_ VPWR VGND _3383_ block[56] round_key[56] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_49_625 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6944_ _2063_ _2397_ _3755_ _2064_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_49_647 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6875_ VPWR VGND VPWR VGND _2155_ _2231_ _2328_ _2327_ _2149_ ZI_sky130_fd_sc_hd__a22oi_2
XFILLER_0_17_500 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5826_ VPWR VGND VGND VPWR _1288_ _3754_ _1287_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_63_105 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_29_393 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5757_ VGND VPWR VGND VPWR _1221_ _0684_ _0609_ _0579_ _0531_ ZI_sky130_fd_sc_hd__and4_2
XFILLER_0_63_149 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_60_81 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_32_525 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8476_ VGND VPWR VPWR VGND clk _0078_ reset_n new_block[35] ZI_sky130_fd_sc_hd__dfrtp_2
X_4708_ VGND VPWR VGND VPWR _0184_ _4134_ _4002_ _0181_ _0183_ ZI_sky130_fd_sc_hd__a211o_2
X_7427_ VGND VPWR _2867_ _0994_ _1126_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5688_ VPWR VGND VPWR VGND _0842_ _1152_ _0924_ _0854_ _1153_ ZI_sky130_fd_sc_hd__or4_2
X_4639_ VGND VPWR VGND VPWR _4114_ _4116_ _3982_ _4021_ _4176_ ZI_sky130_fd_sc_hd__o22a_2
X_7358_ VGND VPWR _2803_ _0994_ _1069_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_580 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6309_ VPWR VGND _1769_ block[18] round_key[18] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7289_ VGND VPWR _2737_ _2735_ _2736_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_113 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_39_146 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_54_127 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_94_274 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_55_628 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_82_447 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_62_193 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_49_16 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_31_580 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_49_49 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_4_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4990_ VPWR VGND VPWR VGND _3946_ _4019_ _4133_ _3913_ _0462_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_81_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_252 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6660_ VPWR VGND _2113_ _2114_ _2060_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5611_ VPWR VGND VPWR VGND _4094_ _1077_ _0366_ _1076_ _1078_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_45_138 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6591_ VGND VPWR VPWR VGND _2044_ _2040_ _2046_ _1277_ _2045_ ZI_sky130_fd_sc_hd__o211a_2
X_5542_ VGND VPWR VGND VPWR _1009_ new_block[106] _1008_ _1003_ _0984_ _0021_ ZI_sky130_fd_sc_hd__o32a_2
X_8330_ VPWR VGND _3687_ _1688_ _1577_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8261_ VGND VPWR _3625_ _3623_ _3624_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5473_ VPWR VGND VPWR VGND _0940_ _0615_ _0939_ _0745_ _0606_ _0941_ ZI_sky130_fd_sc_hd__a221o_2
X_4424_ VGND VPWR _3962_ _3961_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7212_ _2338_ _2661_ _2343_ _2229_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8192_ VGND VPWR VGND VPWR _3563_ _3562_ _3561_ _3558_ ZI_sky130_fd_sc_hd__o21a_2
X_7143_ VPWR VGND VPWR VGND _2361_ _2285_ _2368_ _2169_ _2373_ _2593_ ZI_sky130_fd_sc_hd__a221o_2
X_4355_ VGND VPWR VGND VPWR _3893_ _3892_ _3815_ _3891_ _3890_ ZI_sky130_fd_sc_hd__and4_2
X_7074_ VPWR VGND VGND VPWR _2059_ _2525_ _3776_ ZI_sky130_fd_sc_hd__nor2_2
X_4286_ _3821_ _3824_ _3752_ _3823_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6025_ VGND VPWR _1487_ _1486_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_96_528 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7976_ VPWR VGND VPWR VGND _3309_ _3367_ _3366_ _3328_ _0912_ _3368_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_37_606 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6927_ _2161_ _2380_ _2186_ _2177_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6858_ VPWR VGND _2312_ _2311_ _2310_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_17_330 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5809_ VGND VPWR _1272_ _0794_ _1132_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_107_505 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_91_255 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_64_469 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8528_ VGND VPWR VPWR VGND clk _0130_ reset_n new_block[23] ZI_sky130_fd_sc_hd__dfrtp_2
X_6789_ VPWR VGND VPWR VGND _2211_ _2242_ _2221_ _2185_ _2243_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_91_277 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_44_193 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_91_299 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8459_ VGND VPWR VPWR VGND clk _0061_ reset_n new_block[82] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_388 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_95_594 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_82_233 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_35_160 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_50_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_50_152 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7830_ VGND VPWR VGND VPWR _3234_ _3230_ _3235_ _3028_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_25_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4973_ VPWR VGND _0446_ block[69] round_key[69] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7761_ VGND VPWR _3172_ _2912_ _3171_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7692_ VGND VPWR _3109_ _0381_ _3108_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6712_ _2078_ _2166_ _3754_ _2160_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6643_ VGND VPWR _2097_ _2096_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_46_469 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_73_255 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6574_ VPWR VGND VPWR VGND _1467_ _2028_ _1591_ _1463_ _2029_ ZI_sky130_fd_sc_hd__or4_2
X_8313_ VPWR VGND _3672_ _1234_ _1228_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_14_333 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5525_ VPWR VGND _0993_ round_key[55] new_block[55] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8244_ VGND VPWR VGND VPWR _3610_ _3609_ _3608_ _3605_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_41_163 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5456_ VPWR VGND VGND VPWR _0837_ _0924_ _0622_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_112_585 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4407_ VGND VPWR _3945_ _3815_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_1_271 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8175_ VGND VPWR _3548_ _3461_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5387_ VPWR VGND VGND VPWR _0856_ _0582_ _0698_ ZI_sky130_fd_sc_hd__nand2_2
X_4338_ VPWR VGND VPWR VGND _3809_ _3876_ _3774_ _3814_ ZI_sky130_fd_sc_hd__or3b_2
X_7126_ _2339_ _2576_ _2187_ _2260_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7057_ VGND VPWR VGND VPWR _2508_ _2246_ _2355_ _2205_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_66_80 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4269_ VGND VPWR VPWR VGND sword_ctr_reg\[0\] _3807_ new_block[34] ZI_sky130_fd_sc_hd__and2b_2
X_6008_ VPWR VGND VGND VPWR _1436_ _1470_ _1344_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_69_517 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7959_ VGND VPWR _3352_ _3349_ _3351_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_530 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_103_585 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_62_16 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_43_439 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_102_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6290_ VGND VPWR VPWR VGND _1740_ _1749_ _1724_ _1750_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_51_461 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5310_ VPWR VGND VGND VPWR _0780_ _0582_ _0684_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_87_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5241_ VPWR VGND _0605_ _0711_ _0568_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5172_ VPWR VGND VGND VPWR _0642_ _3914_ _0551_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_78_336 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7813_ VPWR VGND VPWR VGND _3219_ _3159_ _3218_ _3139_ _0794_ _3220_ ZI_sky130_fd_sc_hd__a221o_2
X_7744_ VGND VPWR VPWR VGND _3155_ _1832_ _3157_ _3118_ _3156_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_59_561 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_46_222 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_74_520 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4956_ VPWR VGND VPWR VGND _0417_ _0428_ _0423_ _4167_ _0429_ ZI_sky130_fd_sc_hd__or4_2
X_4887_ VPWR VGND VPWR VGND _0349_ _0360_ _0353_ _0340_ _0361_ ZI_sky130_fd_sc_hd__or4_2
X_7675_ VPWR VGND VPWR VGND _2995_ _2960_ _3093_ _2984_ _0300_ _3094_ ZI_sky130_fd_sc_hd__a221o_2
X_6626_ VGND VPWR VGND VPWR sword_ctr_reg\[0\] new_block[56] sword_ctr_reg\[1\] _2080_
+ ZI_sky130_fd_sc_hd__nand3b_2
XFILLER_0_61_225 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_15_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6557_ VGND VPWR VGND VPWR _1911_ new_block[118] _2012_ _2009_ _1996_ _0033_ ZI_sky130_fd_sc_hd__o32a_2
X_5508_ VPWR VGND VPWR VGND _0731_ _0678_ _0746_ _0635_ _0976_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_30_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6488_ VPWR VGND _1945_ round_key[20] new_block[20] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8227_ VPWR VGND VPWR VGND _3575_ _3490_ _3594_ _3583_ _1689_ _3595_ ZI_sky130_fd_sc_hd__a221o_2
X_5439_ VPWR VGND _0908_ round_key[33] new_block[33] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_100_566 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8158_ VPWR VGND VGND VPWR _3532_ _3521_ _0162_ _3530_ _3531_ _3533_ ZI_sky130_fd_sc_hd__a311o_2
X_7109_ VPWR VGND _2560_ _2497_ _2311_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8089_ VPWR VGND VPWR VGND _3459_ _3367_ _3469_ _3468_ _1684_ _3470_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_96_155 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_96_177 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_96_166 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_52_203 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_65_597 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_80_545 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_20_122 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_103_360 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_21_667 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_88_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_88_634 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_73_48 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4810_ VPWR VGND VGND VPWR _0285_ _0284_ _0283_ _0282_ _4106_ _4046_ ZI_sky130_fd_sc_hd__o2111a_2
X_5790_ VGND VPWR VGND VPWR _0787_ _0619_ _0828_ _1253_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_16_406 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4741_ VGND VPWR VGND VPWR _3976_ _3872_ _3988_ _0217_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_22_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_43_225 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7460_ VGND VPWR _2897_ _1950_ _2896_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4672_ VGND VPWR _0149_ new_block[87] round_key[87] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6411_ VGND VPWR VGND VPWR _1869_ _1444_ _1427_ _1397_ ZI_sky130_fd_sc_hd__o21a_2
X_7391_ VPWR VGND _2833_ _1230_ _0986_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_24_450 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6342_ VPWR VGND VGND VPWR _1800_ _1726_ _1521_ _1474_ _1557_ _1801_ ZI_sky130_fd_sc_hd__a311o_2
XFILLER_0_11_122 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_12_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_98_78 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_11_144 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6273_ VGND VPWR VGND VPWR _1495_ _1371_ _1552_ _1733_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_11_188 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8012_ VGND VPWR VGND VPWR _3399_ _3396_ _3400_ _3339_ ZI_sky130_fd_sc_hd__a21oi_2
X_5224_ VGND VPWR VPWR VGND _0686_ _0693_ _0682_ _0694_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_37_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5155_ VGND VPWR VGND VPWR _0625_ _0585_ _0532_ _0611_ _0624_ ZI_sky130_fd_sc_hd__a211o_2
X_5086_ VPWR VGND VPWR VGND _0556_ new_block[108] _3828_ ZI_sky130_fd_sc_hd__or2_2
XFILLER_0_98_409 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_78_133 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_94_637 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_63_81 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5988_ VPWR VGND VPWR VGND _1429_ _1449_ _1439_ _1423_ _1450_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_93_147 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_93_169 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7727_ VGND VPWR VGND VPWR _2799_ new_block[95] _3141_ _3138_ _2775_ _0074_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_62_501 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4939_ VPWR VGND VGND VPWR _0193_ _0208_ _0412_ ZI_sky130_fd_sc_hd__or2b_2
XFILLER_0_19_277 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_47_597 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7658_ VGND VPWR _3078_ _0369_ _3077_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6609_ VPWR VGND VPWR VGND _2062_ _3764_ _2061_ _3762_ new_block[62] _2063_ ZI_sky130_fd_sc_hd__a221o_2
X_7589_ VGND VPWR _3015_ _3012_ _3014_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_84_125 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_84_114 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_25_225 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_65_361 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_111_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6960_ VGND VPWR _2413_ _0920_ _2412_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_65 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5911_ VPWR VGND VPWR VGND _1372_ _1361_ _1359_ _1337_ _1332_ _1373_ ZI_sky130_fd_sc_hd__a221o_2
X_6891_ VPWR VGND VPWR VGND _2073_ _2330_ _2174_ _2136_ _2344_ ZI_sky130_fd_sc_hd__a22o_2
X_5842_ VPWR VGND VGND VPWR sword_ctr_reg\[0\] sword_ctr_reg\[1\] new_block[115] _1304_
+ ZI_sky130_fd_sc_hd__nor3_2
XFILLER_0_33_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5773_ VGND VPWR _1237_ _1233_ _1236_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_169 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_16_214 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_29_597 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7512_ VGND VPWR _2945_ _1895_ _2944_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4724_ _0185_ _0200_ _3948_ _3934_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8492_ VGND VPWR VPWR VGND clk _0094_ reset_n new_block[51] ZI_sky130_fd_sc_hd__dfrtp_2
X_4655_ VGND VPWR VGND VPWR _4192_ _3857_ _3814_ _3776_ _3804_ ZI_sky130_fd_sc_hd__o211ai_2
X_7443_ VPWR VGND VPWR VGND _2797_ _2881_ _2857_ _2880_ _0295_ _2882_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_71_386 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7374_ VGND VPWR VGND VPWR _2818_ _2817_ _2816_ _2815_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_31_228 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4586_ VPWR VGND VGND VPWR _3964_ _4108_ _4122_ _4123_ ZI_sky130_fd_sc_hd__nor3_2
X_6325_ VGND VPWR VGND VPWR _1784_ _1470_ _1557_ _1782_ _1783_ ZI_sky130_fd_sc_hd__a211o_2
X_6256_ VPWR VGND VPWR VGND _1619_ _1616_ _1438_ _1528_ _1716_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_58_81 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6187_ VPWR VGND VPWR VGND _1645_ _1647_ _1646_ _1644_ _1648_ ZI_sky130_fd_sc_hd__or4_2
X_5207_ VGND VPWR _0677_ _0676_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5138_ VPWR VGND VGND VPWR _3787_ _0608_ _0562_ _0567_ ZI_sky130_fd_sc_hd__nor3b_2
XFILLER_0_98_206 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5069_ VGND VPWR VGND VPWR _0539_ sword_ctr_reg\[0\] new_block[75] sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__and3b_2
XFILLER_0_67_626 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_47_350 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_109_249 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_30_272 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_38_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_100_182 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_445 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_57_125 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_108_260 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_26_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4440_ VPWR VGND VGND VPWR _3978_ _3894_ _3878_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_79_69 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_110_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6110_ VGND VPWR _1572_ _1568_ _1571_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4371_ VPWR VGND VPWR VGND _3889_ _3908_ _3899_ _3867_ _3909_ ZI_sky130_fd_sc_hd__or4_2
X_7090_ VGND VPWR VGND VPWR _2541_ _2223_ _2159_ _2352_ _2540_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_95_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6041_ _1400_ _1503_ _1394_ _1493_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_95_79 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7992_ VGND VPWR VPWR VGND _3380_ _0797_ _3382_ _3265_ _3381_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_44_61 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6943_ VGND VPWR VGND VPWR _2396_ _2196_ _2372_ _2394_ _2395_ ZI_sky130_fd_sc_hd__a211o_2
X_6874_ VGND VPWR _2327_ _2123_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_88_283 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5825_ VGND VPWR VGND VPWR _0538_ _1283_ _1284_ _1285_ _1286_ _1287_ ZI_sky130_fd_sc_hd__o41a_2
XFILLER_0_29_350 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_17_556 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_44_331 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5756_ VPWR VGND VPWR VGND _0828_ _0634_ _1219_ _0713_ _0755_ _1220_ ZI_sky130_fd_sc_hd__a221o_2
X_4707_ VPWR VGND VGND VPWR _4110_ _0183_ _0182_ ZI_sky130_fd_sc_hd__nor2_2
X_5687_ VGND VPWR VGND VPWR _1152_ _0731_ _0740_ _1151_ _0641_ ZI_sky130_fd_sc_hd__a211o_2
X_8475_ VGND VPWR VPWR VGND clk _0077_ reset_n new_block[34] ZI_sky130_fd_sc_hd__dfrtp_2
X_7426_ VPWR VGND _2866_ _1064_ _1068_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4638_ VPWR VGND VGND VPWR _4175_ _3815_ _3920_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_8_61 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_8_94 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7357_ VGND VPWR _2802_ _0914_ _2801_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4569_ VPWR VGND VPWR VGND _4106_ _3865_ _3932_ ZI_sky130_fd_sc_hd__or2_2
X_7288_ VPWR VGND _2736_ _2691_ _1241_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6308_ VGND VPWR VGND VPWR _1768_ _1767_ _1766_ _1758_ ZI_sky130_fd_sc_hd__o21a_2
X_6239_ VGND VPWR VGND VPWR _1699_ _1397_ _1335_ _1697_ _1698_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_39_125 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_39_158 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_67_456 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_67_445 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_55_607 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_94_286 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_49_28 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_81_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_98_581 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_85_220 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_14_53 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_58_467 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5610_ VPWR VGND _1077_ block[43] round_key[43] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6590_ VPWR VGND VGND VPWR _2045_ _2040_ _2044_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_5_225 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5541_ VGND VPWR _1009_ _4103_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_26_353 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_30_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_5_258 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8260_ VGND VPWR _3624_ _0985_ _0998_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_74 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_81_492 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_81_470 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_30_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5472_ VGND VPWR VGND VPWR _0940_ _0638_ _0591_ _0605_ _0582_ ZI_sky130_fd_sc_hd__and4_2
X_7211_ VPWR VGND VPWR VGND _2583_ _2299_ _2355_ _2073_ _2144_ _2660_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_41_389 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8191_ VGND VPWR VGND VPWR _3561_ _3558_ _3562_ _3339_ ZI_sky130_fd_sc_hd__a21oi_2
X_4423_ VGND VPWR _3961_ _3960_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7142_ VPWR VGND VPWR VGND _2589_ _2591_ _2590_ _2588_ _2592_ ZI_sky130_fd_sc_hd__or4_2
X_4354_ VGND VPWR VPWR VGND _3884_ _3883_ _3892_ _3754_ _3843_ ZI_sky130_fd_sc_hd__o211a_2
X_7073_ VPWR VGND VPWR VGND _2457_ _2523_ _2522_ _2521_ _2524_ ZI_sky130_fd_sc_hd__or4_2
X_6024_ VPWR VGND VPWR VGND _1393_ _1388_ _1288_ _1391_ _1486_ ZI_sky130_fd_sc_hd__or4_2
X_4285_ VPWR VGND VPWR VGND _3823_ new_block[103] _3822_ ZI_sky130_fd_sc_hd__or2_2
X_7975_ VGND VPWR _3367_ _0161_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6926_ VPWR VGND _2149_ _2379_ _2204_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_76_220 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6857_ VPWR VGND _2311_ new_block[127] round_key[127] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5808_ VGND VPWR _1271_ _0802_ _1188_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6788_ VPWR VGND VPWR VGND _2226_ _2241_ _2232_ _2224_ _2242_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_107_517 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8527_ VGND VPWR VPWR VGND clk _0129_ reset_n new_block[22] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_651 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_51_109 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5739_ VGND VPWR VGND VPWR _1203_ _0765_ _0662_ _1200_ _1202_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_44_183 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_91_289 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_60_610 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8458_ VGND VPWR VPWR VGND clk _0060_ reset_n new_block[81] ZI_sky130_fd_sc_hd__dfrtp_2
X_7409_ VGND VPWR _2850_ _0808_ _2849_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8389_ VPWR VGND VPWR VGND _3521_ _4093_ _3740_ _0169_ _1680_ _3741_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_35_19 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_59_209 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_82_245 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_42_109 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_51_654 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_50_164 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_50_197 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4972_ VGND VPWR VPWR VGND _0442_ _0433_ _0445_ _0444_ _0443_ ZI_sky130_fd_sc_hd__o211a_2
X_7760_ VPWR VGND _3171_ _1818_ _1576_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_19_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7691_ VGND VPWR _3108_ _4072_ _4076_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6711_ VPWR VGND _2150_ _2165_ _2164_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_73_201 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_58_253 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_41_40 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6642_ VPWR VGND VGND VPWR _2095_ _2096_ _2084_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_73_267 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6573_ VPWR VGND VPWR VGND _1419_ _1778_ _1341_ _1471_ _2028_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_6_578 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8312_ VGND VPWR _3671_ _1272_ _3670_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5524_ VPWR VGND _0992_ round_key[50] new_block[50] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8243_ VGND VPWR VGND VPWR _3608_ _3605_ _3609_ _4085_ ZI_sky130_fd_sc_hd__a21oi_2
X_5455_ VGND VPWR _0923_ _0688_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8174_ VPWR VGND VPWR VGND _3459_ _3490_ _3546_ _3468_ _1688_ _3547_ ZI_sky130_fd_sc_hd__a221o_2
X_4406_ VGND VPWR VGND VPWR _3939_ _3938_ _3943_ _3944_ ZI_sky130_fd_sc_hd__a21o_2
X_7125_ VPWR VGND VPWR VGND _2097_ _2184_ _2112_ _2255_ _2575_ ZI_sky130_fd_sc_hd__a22o_2
X_5386_ VGND VPWR VGND VPWR _0855_ _0596_ _0854_ _0736_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_5_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4337_ VPWR VGND VGND VPWR _3874_ _3875_ _3854_ ZI_sky130_fd_sc_hd__nor2_2
X_7056_ VPWR VGND _2174_ _2507_ _2259_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_4268_ sword_ctr_reg\[1\] _3806_ sword_ctr_reg\[0\] new_block[2] VPWR VGND VPWR VGND
+ ZI_sky130_fd_sc_hd__and3_2
X_6007_ VGND VPWR VGND VPWR _1469_ _1464_ _1341_ _1467_ _1468_ ZI_sky130_fd_sc_hd__a211o_2
X_4199_ VPWR VGND VGND VPWR _3748_ dec_ctrl_reg\[0\] next ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_96_326 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_69_529 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7958_ VGND VPWR _3351_ _4069_ _3350_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7889_ VGND VPWR _3288_ _0489_ _2312_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6909_ VPWR VGND VPWR VGND _2361_ _2201_ _2281_ _2169_ _2176_ _2362_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_77_584 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_59_Left_172 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_37_437 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_64_223 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_33_643 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_103_542 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_20_359 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_103_597 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_181 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_99_164 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_77_Left_190 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_68_573 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_55_201 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_15_109 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_51_473 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5240_ VGND VPWR _0710_ _0709_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_18_Right_18 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5171_ VPWR VGND VGND VPWR _0640_ _0641_ _0637_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_78_348 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7812_ VGND VPWR _3219_ _3149_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_27_Right_27 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7743_ VPWR VGND VGND VPWR _3156_ _1832_ _3155_ ZI_sky130_fd_sc_hd__nand2_2
X_4955_ VPWR VGND VPWR VGND _4108_ _0427_ _0424_ _3889_ _0428_ ZI_sky130_fd_sc_hd__or4_2
X_4886_ VPWR VGND VPWR VGND _0358_ _0359_ _0360_ _0354_ _0355_ ZI_sky130_fd_sc_hd__or4b_2
X_7674_ VPWR VGND _3093_ block[91] round_key[91] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6625_ VGND VPWR VGND VPWR new_block[24] sword_ctr_reg\[0\] _2079_ sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__nand3_2
X_6556_ VPWR VGND VPWR VGND _1281_ _1909_ _2011_ _1959_ _2010_ _2012_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_15_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5507_ VGND VPWR _0975_ _0939_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_42_473 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_30_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8226_ VPWR VGND _3594_ block[78] round_key[78] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_112_361 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6487_ VPWR VGND _1944_ _1891_ _1820_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_36_Right_36 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5438_ VPWR VGND _0907_ round_key[38] new_block[38] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8157_ VPWR VGND VGND VPWR _1683_ _3532_ _4089_ ZI_sky130_fd_sc_hd__nor2_2
X_5369_ VPWR VGND VGND VPWR _0724_ _0838_ _0837_ ZI_sky130_fd_sc_hd__nor2_2
X_7108_ VGND VPWR _2559_ _2556_ _2558_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_578 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_100_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8088_ VPWR VGND _3469_ block[97] round_key[97] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7039_ VPWR VGND _2491_ _2490_ _2409_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_93_90 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_108_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_52_226 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_108_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_92_384 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_21_613 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_54_Right_54 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Right_63 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_88_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_87_123 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4740_ VPWR VGND VGND VPWR _4181_ _4116_ _3984_ _4114_ _0216_ _0215_ ZI_sky130_fd_sc_hd__o221a_2
XFILLER_0_56_565 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_56_543 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4671_ VPWR VGND _0148_ _0147_ _4068_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6410_ VPWR VGND VPWR VGND _1867_ _1534_ _1626_ _1375_ _1546_ _1868_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_43_237 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7390_ VGND VPWR VGND VPWR _2800_ new_block[67] _2832_ _2830_ _0294_ _0046_ ZI_sky130_fd_sc_hd__o32a_2
X_6341_ VPWR VGND VPWR VGND _1534_ _1629_ _1430_ _1636_ _1800_ ZI_sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_72_Right_72 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_71_579 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6272_ VGND VPWR VGND VPWR _1732_ _1639_ _1471_ _1606_ _1731_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_11_134 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_12_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8011_ VGND VPWR _3399_ _0987_ _3398_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5223_ VGND VPWR VGND VPWR _0693_ _0677_ _0689_ _0692_ _0690_ _0688_ ZI_sky130_fd_sc_hd__a32o_2
X_5154_ VPWR VGND VPWR VGND _0623_ _0607_ _0619_ _0613_ _0616_ _0624_ ZI_sky130_fd_sc_hd__a221o_2
X_5085_ VGND VPWR VGND VPWR _0555_ _0552_ _3764_ _0553_ _0554_ ZI_sky130_fd_sc_hd__a211o_2
XPHY_EDGE_ROW_81_Right_81 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_63_93 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_19_212 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5987_ VPWR VGND VPWR VGND _1448_ _1332_ _1443_ _1440_ _1421_ _1449_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_47_532 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_93_126 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_19_245 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4938_ VGND VPWR VGND VPWR _0218_ _4030_ _0406_ _0408_ _0411_ _0410_ ZI_sky130_fd_sc_hd__a2111o_2
X_7726_ VPWR VGND VPWR VGND _2995_ _3140_ _0162_ _3139_ _4061_ _3141_ ZI_sky130_fd_sc_hd__a221o_2
X_4869_ VGND VPWR VGND VPWR _0343_ _0218_ _3946_ _0341_ _0342_ ZI_sky130_fd_sc_hd__a211o_2
X_7657_ VGND VPWR _3077_ _0232_ _3076_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_248 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_90_Right_90 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6608_ sword_ctr_reg\[1\] _2062_ sword_ctr_reg\[0\] new_block[30] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
X_7588_ VGND VPWR _3014_ _2487_ _3013_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6539_ VPWR VGND VPWR VGND _1983_ _1994_ _1986_ _1976_ _1995_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_30_421 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8209_ VGND VPWR _3578_ _3086_ _3577_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_69_178 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_69_156 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_84_137 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_65_373 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_80_365 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_68_16 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_21_443 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_111_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_108_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5910_ VPWR VGND VGND VPWR _1371_ _1372_ _1366_ ZI_sky130_fd_sc_hd__nor2_2
X_6890_ VGND VPWR _2343_ _2127_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5841_ VPWR VGND VGND VPWR sword_ctr_reg\[0\] new_block[51] _1303_ ZI_sky130_fd_sc_hd__or2b_2
X_5772_ VGND VPWR _1236_ _1234_ _1235_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8491_ VGND VPWR VPWR VGND clk _0093_ reset_n new_block[50] ZI_sky130_fd_sc_hd__dfrtp_2
X_7511_ VPWR VGND _2944_ _2915_ _1565_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4723_ VGND VPWR VGND VPWR _4143_ _3804_ _0196_ _0197_ _0199_ _0198_ ZI_sky130_fd_sc_hd__a2111o_2
X_7442_ VPWR VGND _2881_ block[39] round_key[39] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4654_ _3804_ _4191_ _3894_ _3950_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7373_ VGND VPWR VGND VPWR _2816_ _2815_ _2817_ _2642_ ZI_sky130_fd_sc_hd__a21oi_2
X_4585_ VPWR VGND VPWR VGND _4120_ _4121_ _4122_ _4113_ _4118_ ZI_sky130_fd_sc_hd__or4b_2
X_6324_ VGND VPWR VGND VPWR _1501_ _1522_ _1487_ _1462_ _1783_ ZI_sky130_fd_sc_hd__a2bb2o_2
X_6255_ VPWR VGND VPWR VGND _1712_ _1714_ _1713_ _1503_ _1715_ ZI_sky130_fd_sc_hd__or4_2
X_5206_ _0643_ _0676_ _0642_ _0608_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6186_ _1455_ _1647_ _1394_ _1530_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5137_ VGND VPWR _0607_ _0606_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_98_218 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5068_ VGND VPWR _0538_ _3788_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Right_0 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7709_ VGND VPWR _3125_ _0384_ _0482_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_660 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_50_516 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_100_161 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_89_207 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_72_107 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_81_630 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_65_181 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_108_272 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4370_ VGND VPWR VGND VPWR _3907_ _3795_ _3900_ _3903_ _3908_ ZI_sky130_fd_sc_hd__a31o_2
XPHY_EDGE_ROW_13_Left_126 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6040_ VGND VPWR VGND VPWR _1502_ _1434_ _1501_ _1443_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_28_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7991_ VPWR VGND VGND VPWR _3381_ _0797_ _3380_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_44_40 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6942_ VPWR VGND VPWR VGND _2279_ _2368_ _2260_ _2236_ _2395_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_44_73 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6873_ VPWR VGND VPWR VGND _2203_ _2326_ _2166_ _2225_ ZI_sky130_fd_sc_hd__or3b_2
XPHY_EDGE_ROW_22_Left_135 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5824_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[112] sword_ctr_reg\[0\] _1286_
+ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_48_148 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5755_ VPWR VGND _0620_ _1219_ _0827_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_106_209 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_56_181 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_97_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_71_140 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4706_ VPWR VGND VGND VPWR _0182_ _3804_ _3881_ ZI_sky130_fd_sc_hd__nand2_2
X_8474_ VGND VPWR VPWR VGND clk _0076_ reset_n new_block[33] ZI_sky130_fd_sc_hd__dfrtp_2
X_5686_ VPWR VGND VPWR VGND _0678_ _0658_ _0627_ _0666_ _1151_ ZI_sky130_fd_sc_hd__a22o_2
X_7425_ VGND VPWR _2865_ _2863_ _2864_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4637_ VPWR VGND VPWR VGND _4174_ _4167_ _4173_ ZI_sky130_fd_sc_hd__or2_2
X_7356_ VGND VPWR _2801_ _0801_ _0998_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4568_ VPWR VGND VGND VPWR _4105_ _3881_ _3925_ ZI_sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_31_Left_144 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4499_ VGND VPWR VGND VPWR _4022_ _3862_ _4037_ _4036_ ZI_sky130_fd_sc_hd__a21oi_2
X_7287_ VGND VPWR _2735_ _2565_ _2734_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6307_ VGND VPWR VGND VPWR _1766_ _1758_ _1767_ _1001_ ZI_sky130_fd_sc_hd__a21oi_2
X_6238_ VPWR VGND VGND VPWR _1547_ _1698_ _1366_ ZI_sky130_fd_sc_hd__nor2_2
X_6169_ VGND VPWR VGND VPWR _1630_ _1395_ _1531_ _1397_ ZI_sky130_fd_sc_hd__o21a_2
XPHY_EDGE_ROW_40_Left_153 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_39_104 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_63_641 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_23_505 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_62_173 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_81_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_14_98 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5540_ VGND VPWR VGND VPWR _1007_ _4094_ _1004_ _1005_ _1008_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_30_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5471_ VPWR VGND VGND VPWR _0655_ _0939_ _0617_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_30_97 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7210_ VGND VPWR VGND VPWR _2659_ _2159_ _2216_ _2369_ _2450_ ZI_sky130_fd_sc_hd__a211o_2
X_4422_ VPWR VGND VPWR VGND _3901_ _3960_ _3830_ _3863_ ZI_sky130_fd_sc_hd__or3b_2
X_8190_ VGND VPWR _3561_ _3083_ _3560_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_40 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7141_ VGND VPWR VGND VPWR _2591_ _2300_ _2256_ _2190_ ZI_sky130_fd_sc_hd__o21a_2
X_4353_ VGND VPWR _3891_ _3863_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7072_ _2166_ _2523_ _2186_ _2267_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_4284_ VPWR VGND VPWR VGND _3822_ sword_ctr_reg\[0\] sword_ctr_reg\[1\] ZI_sky130_fd_sc_hd__or2_2
X_6023_ VPWR VGND VPWR VGND _1463_ _1484_ _1469_ _1458_ _1485_ ZI_sky130_fd_sc_hd__or4_2
X_7974_ VPWR VGND _3366_ block[86] round_key[86] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_12_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_49_424 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6925_ _2162_ _2378_ _2070_ _2175_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6856_ VPWR VGND _2310_ new_block[125] round_key[125] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5807_ VGND VPWR _1270_ _1228_ _1269_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6787_ VGND VPWR VGND VPWR _2194_ _2233_ _2234_ _2238_ _2241_ _2240_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_64_438 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8526_ VGND VPWR VPWR VGND clk _0128_ reset_n new_block[21] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_663 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_107_529 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5738_ VPWR VGND VPWR VGND _1201_ _0704_ _0736_ _0669_ _0975_ _1202_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_60_622 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5669_ VPWR VGND _1135_ _0988_ _0902_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8457_ VGND VPWR VPWR VGND clk _0059_ reset_n new_block[80] ZI_sky130_fd_sc_hd__dfrtp_2
X_7408_ VPWR VGND _2849_ _1137_ _0805_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8388_ VPWR VGND _3740_ block[30] round_key[30] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7339_ VGND VPWR _2786_ _0161_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_102_289 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_55_449 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_51_633 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_92_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4971_ VGND VPWR _0444_ _0365_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7690_ VGND VPWR _3107_ _0239_ _0373_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_585 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6710_ VPWR VGND VPWR VGND _2103_ _2163_ _2161_ _2162_ _2164_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_58_265 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_18_118 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6641_ VGND VPWR VGND VPWR _2094_ _2089_ _2095_ _3850_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_58_287 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_27_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_41_52 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6572_ VPWR VGND VPWR VGND _1982_ _2026_ _2025_ _1631_ _2027_ ZI_sky130_fd_sc_hd__or4_2
X_8311_ VPWR VGND _3670_ _0800_ _0795_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_41_96 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5523_ VGND VPWR _0991_ _0987_ _0990_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5454_ VGND VPWR VGND VPWR _4104_ new_block[105] _0922_ _0917_ _0899_ _0020_ ZI_sky130_fd_sc_hd__o32a_2
X_8242_ VGND VPWR _3608_ _3606_ _3607_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5385_ VGND VPWR VGND VPWR _0854_ _0569_ _0643_ _0642_ _0579_ ZI_sky130_fd_sc_hd__and4_2
X_4405_ VPWR VGND VGND VPWR _3942_ _3943_ _3941_ ZI_sky130_fd_sc_hd__nor2_2
X_8173_ VPWR VGND _3546_ block[73] round_key[73] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7124_ VPWR VGND VPWR VGND _2511_ _2573_ _2570_ _2359_ _2574_ ZI_sky130_fd_sc_hd__or4_2
X_4336_ VPWR VGND VPWR VGND _3838_ _3847_ _3824_ _3831_ _3874_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_10_596 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7055_ VPWR VGND VPWR VGND _2505_ _2338_ _2155_ _2174_ _2222_ _2506_ ZI_sky130_fd_sc_hd__a221o_2
X_4267_ VGND VPWR VGND VPWR _3805_ sword_ctr_reg\[0\] new_block[66] sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__and3b_2
X_6006_ VGND VPWR VGND VPWR _1468_ _1340_ _1351_ _1345_ ZI_sky130_fd_sc_hd__o21a_2
X_7957_ VPWR VGND _3350_ _0367_ _0305_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7888_ VGND VPWR VGND VPWR _3240_ new_block[46] _3287_ _3285_ _1227_ _0089_ ZI_sky130_fd_sc_hd__o32a_2
X_6908_ VGND VPWR VGND VPWR _2361_ _2175_ _2139_ _2129_ _2117_ ZI_sky130_fd_sc_hd__and4_2
XFILLER_0_37_449 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6839_ VPWR VGND VPWR VGND _2284_ _2292_ _2287_ _2283_ _2293_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_107_337 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_33_611 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_33_655 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8509_ VGND VPWR VPWR VGND clk _0111_ reset_n new_block[4] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_305 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_103_554 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_1_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_99_176 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_83_544 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_68_585 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_70_205 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_23_154 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_87_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_23_187 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_51_485 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5170_ VPWR VGND VGND VPWR _0640_ _0545_ _0639_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_36_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_36_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7811_ VPWR VGND _3218_ block[7] round_key[7] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7742_ VGND VPWR _3155_ _2929_ _3154_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4954_ VPWR VGND VGND VPWR _0426_ _0425_ _4008_ _3934_ _4012_ _0427_ ZI_sky130_fd_sc_hd__a311o_2
XFILLER_0_19_449 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4885_ VGND VPWR VGND VPWR _4106_ _0177_ _3920_ _3976_ _3932_ _0359_ ZI_sky130_fd_sc_hd__o32a_2
X_7673_ VGND VPWR VGND VPWR _3092_ _3091_ _3090_ _3089_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_15_611 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6624_ VGND VPWR VGND VPWR _2078_ _4097_ _2074_ _2075_ _2076_ _2077_ ZI_sky130_fd_sc_hd__a41o_2
XFILLER_0_61_216 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_61_205 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_6_365 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6555_ VPWR VGND _2011_ new_block[118] round_key[118] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5506_ VGND VPWR VGND VPWR _0974_ _0778_ _0596_ _0880_ _0973_ ZI_sky130_fd_sc_hd__a211o_2
XPHY_EDGE_ROW_5_Left_118 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6486_ VGND VPWR VPWR VGND _1937_ _1942_ _1930_ _1943_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_30_636 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8225_ VGND VPWR VGND VPWR _3593_ _3592_ _3591_ _3590_ ZI_sky130_fd_sc_hd__o21a_2
X_5437_ VGND VPWR _0906_ _0901_ _0905_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5368_ VPWR VGND VGND VPWR _0837_ _0532_ _0579_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_77_81 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8156_ VPWR VGND VPWR VGND _3531_ round_key[103] block[103] ZI_sky130_fd_sc_hd__or2_2
X_7107_ VPWR VGND _2558_ _2557_ _4087_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5299_ VPWR VGND VPWR VGND _0766_ _0768_ _0769_ _0762_ _0764_ ZI_sky130_fd_sc_hd__or4b_2
X_8087_ VGND VPWR _3468_ _2702_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4319_ VGND VPWR _3857_ _3856_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7038_ VPWR VGND _2490_ _2048_ _1770_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_108_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_9_192 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_108_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_80_503 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_52_249 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4670_ VPWR VGND _0147_ round_key[64] new_block[64] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_56_577 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_3_313 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6340_ VPWR VGND VPWR VGND _1795_ _1798_ _1796_ _1793_ _1799_ ZI_sky130_fd_sc_hd__or4_2
X_6271_ VPWR VGND VPWR VGND _1443_ _1616_ _1464_ _1511_ _1731_ ZI_sky130_fd_sc_hd__a22o_2
X_8010_ VGND VPWR _3398_ _0994_ _3397_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5222_ VGND VPWR _0692_ _0691_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5153_ VPWR VGND VGND VPWR _0622_ _0623_ _0621_ ZI_sky130_fd_sc_hd__nor2_2
X_5084_ sword_ctr_reg\[1\] _0554_ sword_ctr_reg\[0\] new_block[12] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_2_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_2_75 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5986_ VPWR VGND VGND VPWR _1447_ _1448_ _1445_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_47_500 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_19_257 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4937_ VPWR VGND VGND VPWR _0410_ _3957_ _0409_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_47_544 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7725_ VPWR VGND _3140_ block[95] round_key[95] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_7_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4868_ VGND VPWR VGND VPWR _4178_ _4025_ _0342_ _3962_ ZI_sky130_fd_sc_hd__a21oi_2
X_7656_ VPWR VGND _3076_ _0142_ _4063_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6607_ VPWR VGND VGND VPWR new_block[94] sword_ctr_reg\[0\] _2061_ ZI_sky130_fd_sc_hd__or2b_2
XFILLER_0_62_558 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7587_ VPWR VGND _3013_ _2739_ _2630_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4799_ VGND VPWR VGND VPWR _0274_ _0267_ _3949_ _0271_ _0273_ ZI_sky130_fd_sc_hd__a211o_2
X_6538_ VPWR VGND VPWR VGND _1990_ _1993_ _1992_ _1628_ _1994_ ZI_sky130_fd_sc_hd__or4_2
X_6469_ VGND VPWR VGND VPWR _1547_ _1371_ _1926_ _1405_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_30_488 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_112_181 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8208_ VGND VPWR _3577_ _4074_ _3123_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8139_ VGND VPWR _3515_ _3512_ _3514_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_365 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_102_Right_102 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_97_444 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_69_113 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_97_499 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_53_569 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_80_377 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_0_305 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_84_16 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5840_ VGND VPWR VGND VPWR new_block[19] sword_ctr_reg\[0\] _1302_ sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__nand3_2
X_5771_ VPWR VGND _1235_ _1138_ _0801_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_75_138 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8490_ VGND VPWR VPWR VGND clk _0092_ reset_n new_block[49] ZI_sky130_fd_sc_hd__dfrtp_2
X_7510_ VGND VPWR _2943_ _2938_ _2942_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4722_ VPWR VGND VGND VPWR _4121_ _0198_ _3998_ ZI_sky130_fd_sc_hd__nor2_2
X_7441_ VGND VPWR _2880_ _2702_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_44_525 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_44_558 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4653_ VPWR VGND VPWR VGND _4133_ _4041_ _4189_ _3997_ _4190_ ZI_sky130_fd_sc_hd__a22o_2
X_7372_ VGND VPWR _2816_ _0796_ _0909_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4584_ VPWR VGND VPWR VGND _4121_ _3877_ _3920_ ZI_sky130_fd_sc_hd__or2_2
X_6323_ VPWR VGND VGND VPWR _1552_ _1782_ _1475_ ZI_sky130_fd_sc_hd__nor2_2
X_6254_ VPWR VGND VPWR VGND _1426_ _1471_ _1354_ _1456_ _1714_ ZI_sky130_fd_sc_hd__a22o_2
X_5205_ VPWR VGND VGND VPWR _0649_ _0675_ _0532_ ZI_sky130_fd_sc_hd__nor2_2
X_6185_ VGND VPWR VGND VPWR _1646_ _1397_ _1588_ _1421_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_42_3 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_95_Left_208 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5136_ VPWR VGND _0581_ _0606_ _0605_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5067_ VGND VPWR VGND VPWR _3788_ _0533_ _0534_ _0535_ _0537_ _0536_ ZI_sky130_fd_sc_hd__o41ai_2
X_5969_ VPWR VGND VPWR VGND _1431_ _1430_ ZI_sky130_fd_sc_hd__inv_2
X_7708_ VGND VPWR _3124_ _0440_ _3123_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_193 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7639_ VGND VPWR VGND VPWR _3061_ _3060_ _3059_ _0148_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_50_528 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_50_539 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_101_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_100_173 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_97_241 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_97_296 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_70_29 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_81_642 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_108_284 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_80_130 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_79_16 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_80_163 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_21_230 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_95_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_28_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7990_ VGND VPWR _3380_ _2862_ _3379_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_44_52 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6941_ VPWR VGND VPWR VGND _2393_ _2096_ _2260_ _2190_ _2102_ _2394_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_49_617 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6872_ VPWR VGND VPWR VGND _2297_ _2231_ _2302_ _2265_ _2325_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_76_414 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5823_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] _1285_ new_block[80] ZI_sky130_fd_sc_hd__and2b_2
XFILLER_0_8_235 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5754_ VGND VPWR VGND VPWR _0770_ _0633_ _0788_ _0672_ _1218_ _0749_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_60_73 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_71_152 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4705_ VPWR VGND VGND VPWR _3987_ _0181_ _3882_ ZI_sky130_fd_sc_hd__nor2_2
X_5685_ VPWR VGND VPWR VGND _1149_ _0748_ _1148_ _0923_ _1081_ _1150_ ZI_sky130_fd_sc_hd__a221o_2
X_8473_ VGND VPWR VPWR VGND clk _0075_ reset_n new_block[32] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_56_193 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_8_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7424_ VGND VPWR _2864_ _0795_ _1133_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4636_ VPWR VGND VPWR VGND _4170_ _4172_ _4171_ _4169_ _4173_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_71_196 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7355_ VGND VPWR VGND VPWR _2800_ new_block[64] _2798_ _2794_ _4060_ _0043_ ZI_sky130_fd_sc_hd__o32a_2
X_6306_ VGND VPWR _1766_ _1761_ _1765_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4567_ VGND VPWR VGND VPWR _4104_ new_block[96] _4102_ _4091_ _4060_ _0011_ ZI_sky130_fd_sc_hd__o32a_2
X_7286_ VPWR VGND _2734_ _2646_ _2311_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_110_460 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4498_ VGND VPWR _4036_ _4035_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6237_ VPWR VGND VPWR VGND _1471_ _1531_ _1394_ _1379_ _1697_ ZI_sky130_fd_sc_hd__a22o_2
X_6168_ VPWR VGND VGND VPWR _1495_ _1629_ _1366_ ZI_sky130_fd_sc_hd__nor2_2
X_5119_ VGND VPWR _0589_ _0588_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6099_ VPWR VGND VPWR VGND _1517_ _1560_ _1541_ _1505_ _1561_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_79_230 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_94_222 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_62_141 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_105_221 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_62_185 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_81_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_105_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_58_458 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_14_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_30_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5470_ VGND VPWR VGND VPWR _0938_ _0859_ _0662_ _0935_ _0937_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_100_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4421_ VGND VPWR VGND VPWR _3802_ _3793_ _3776_ _3959_ ZI_sky130_fd_sc_hd__a21o_2
X_7140_ VPWR VGND VPWR VGND _2115_ _2279_ _2135_ _2235_ _2590_ ZI_sky130_fd_sc_hd__a22o_2
X_4352_ VGND VPWR _3890_ _3846_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7071_ VGND VPWR VGND VPWR _2522_ _2267_ _2201_ _2106_ ZI_sky130_fd_sc_hd__o21a_2
X_4283_ VGND VPWR VGND VPWR _3821_ _3818_ _3764_ _3819_ _3820_ ZI_sky130_fd_sc_hd__a211o_2
X_6022_ VPWR VGND VPWR VGND _1481_ _1483_ _1482_ _1477_ _1484_ ZI_sky130_fd_sc_hd__or4_2
X_7973_ VGND VPWR VPWR VGND _3363_ _3358_ _3365_ _3265_ _3364_ ZI_sky130_fd_sc_hd__o211a_2
X_6924_ VPWR VGND VPWR VGND _2371_ _2376_ _2375_ _2367_ _2377_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_49_436 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6855_ VPWR VGND _2309_ new_block[126] round_key[126] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_71_83 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5806_ VGND VPWR _1269_ _0805_ _0907_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_555 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_91_225 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6786_ VPWR VGND _2169_ _2240_ _2239_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_8525_ VGND VPWR VPWR VGND clk _0127_ reset_n new_block[20] ZI_sky130_fd_sc_hd__dfrtp_2
X_5737_ VGND VPWR VGND VPWR _1201_ _0695_ _0661_ _0706_ ZI_sky130_fd_sc_hd__o21a_2
X_8456_ VGND VPWR VPWR VGND clk _0058_ reset_n new_block[79] ZI_sky130_fd_sc_hd__dfrtp_2
X_7407_ VPWR VGND _2848_ _1135_ _0811_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5668_ VGND VPWR _1134_ _1131_ _1133_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5599_ VPWR VGND _1066_ _1065_ _0807_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8387_ VPWR VGND VGND VPWR _3738_ _3739_ _3737_ ZI_sky130_fd_sc_hd__nor2_2
X_4619_ VPWR VGND VPWR VGND _4152_ _4155_ _4156_ _3944_ _4150_ ZI_sky130_fd_sc_hd__or4b_2
X_7338_ VPWR VGND _2785_ block[127] round_key[127] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7269_ VGND VPWR VGND VPWR _2717_ _2716_ _2343_ _2590_ _2438_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_67_233 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_50_122 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_23_358 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_50_188 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4970_ VPWR VGND VGND VPWR _0443_ _0433_ _0442_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_46_417 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6640_ VGND VPWR VGND VPWR _0538_ _2090_ _2091_ _2092_ _2094_ _2093_ ZI_sky130_fd_sc_hd__o41ai_2
X_6571_ VPWR VGND VPWR VGND _1792_ _1881_ _2026_ _1429_ _1715_ ZI_sky130_fd_sc_hd__or4b_2
XFILLER_0_27_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_73_247 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5522_ VGND VPWR _0990_ _0908_ _0989_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8310_ VGND VPWR _3669_ _0913_ _1126_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_42_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5453_ VGND VPWR VGND VPWR _0921_ _4094_ _0918_ _0919_ _0922_ ZI_sky130_fd_sc_hd__a31o_2
X_8241_ VGND VPWR _3607_ _0796_ _1192_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_533 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5384_ VGND VPWR VGND VPWR _0851_ _0570_ _0852_ _0853_ ZI_sky130_fd_sc_hd__a21o_2
X_4404_ VGND VPWR VPWR VGND _3878_ _3929_ _3857_ _3942_ ZI_sky130_fd_sc_hd__or3_2
X_8172_ VGND VPWR VPWR VGND _3543_ _3542_ _3545_ _3448_ _3544_ ZI_sky130_fd_sc_hd__o211a_2
X_7123_ VPWR VGND VPWR VGND _2572_ _2118_ _2571_ _2339_ _2198_ _2573_ ZI_sky130_fd_sc_hd__a221o_2
X_4335_ VPWR VGND VGND VPWR _3872_ _3873_ _3870_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_5_97 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7054_ VPWR VGND VPWR VGND _2214_ _2336_ _2120_ _2073_ _2505_ ZI_sky130_fd_sc_hd__a22o_2
X_4266_ VGND VPWR _3804_ _3803_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6005_ VPWR VGND VGND VPWR _1466_ _1467_ _1371_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_49_233 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7956_ VPWR VGND _3349_ _0377_ _0233_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_82_93 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7887_ VPWR VGND VPWR VGND _3219_ _3257_ _3286_ _3237_ _0800_ _3287_ ZI_sky130_fd_sc_hd__a221o_2
X_6907_ VPWR VGND _2114_ _2360_ _2227_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_18_620 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6838_ VPWR VGND VPWR VGND _2289_ _2291_ _2290_ _2288_ _2292_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_9_363 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6769_ VPWR VGND VGND VPWR _2146_ _2223_ _2084_ ZI_sky130_fd_sc_hd__nor2_2
X_8508_ VGND VPWR VPWR VGND clk _0110_ reset_n new_block[3] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_185 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_33_667 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8439_ VGND VPWR VPWR VGND clk _0041_ reset_n new_block[126] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_68_542 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_83_501 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_24_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_51_497 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_87_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_36_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7810_ VGND VPWR VPWR VGND _3215_ _3212_ _3217_ _3118_ _3216_ ZI_sky130_fd_sc_hd__o211a_2
X_7741_ VGND VPWR _3154_ _1828_ _2919_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4953_ VGND VPWR VGND VPWR _3962_ _3896_ _0426_ _3974_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_52_74 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7672_ VGND VPWR VGND VPWR _3090_ _3089_ _3091_ _3028_ ZI_sky130_fd_sc_hd__a21oi_2
X_4884_ VGND VPWR VGND VPWR _0266_ _4008_ _0356_ _0357_ _0358_ _0192_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_52_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6623_ VPWR VGND VGND VPWR sword_ctr_reg\[0\] sword_ctr_reg\[1\] new_block[121] _2077_
+ ZI_sky130_fd_sc_hd__nor3_2
X_6554_ VPWR VGND _2010_ block[22] round_key[22] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_6_377 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_14_111 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6485_ VPWR VGND VPWR VGND _1730_ _1941_ _1732_ _1651_ _1942_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_6_399 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5505_ VGND VPWR VGND VPWR _0973_ _0741_ _0626_ _0643_ ZI_sky130_fd_sc_hd__and3b_2
X_5436_ VPWR VGND _0905_ _0904_ _0902_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8224_ VGND VPWR VGND VPWR _3591_ _3590_ _3592_ _4085_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_72_3 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8155_ VPWR VGND VGND VPWR _3530_ round_key[103] block[103] ZI_sky130_fd_sc_hd__nand2_2
X_5367_ VPWR VGND VPWR VGND _0705_ _0648_ _0836_ _0675_ _0835_ ZI_sky130_fd_sc_hd__or4b_2
X_8086_ VGND VPWR VPWR VGND _3465_ _3463_ _3467_ _3448_ _3466_ ZI_sky130_fd_sc_hd__o211a_2
X_5298_ VGND VPWR VGND VPWR _0589_ _0767_ _0768_ _0688_ _0705_ _0645_ ZI_sky130_fd_sc_hd__a32oi_2
XFILLER_0_77_93 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7106_ VPWR VGND _2557_ _0523_ _0447_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4318_ VPWR VGND VPWR VGND _3856_ _3832_ _3793_ ZI_sky130_fd_sc_hd__or2_2
X_7037_ VGND VPWR _2489_ _2486_ _2488_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4249_ VGND VPWR _3787_ _3773_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7939_ VPWR VGND _3333_ _0374_ _0309_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_106_Left_219 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_77_383 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_108_625 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_18_472 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_107_113 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_87_169 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_83_320 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_56_589 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_98_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_12_604 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6270_ VGND VPWR VGND VPWR _1550_ _1534_ _1729_ _1730_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_11_169 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5221_ VPWR VGND _0598_ _0691_ _0591_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5152_ VPWR VGND VGND VPWR _0622_ _0582_ _0583_ ZI_sky130_fd_sc_hd__nand2_2
X_5083_ VGND VPWR VPWR VGND sword_ctr_reg\[0\] _0553_ new_block[44] ZI_sky130_fd_sc_hd__and2b_2
XFILLER_0_79_604 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_63_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_66_309 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7724_ VGND VPWR _3139_ _2702_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5985_ VGND VPWR _1447_ _1446_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_19_225 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4936_ VGND VPWR VGND VPWR _4115_ _3932_ _3906_ _0409_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_47_556 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_19_269 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4867_ VPWR VGND VGND VPWR _0182_ _0341_ _3906_ ZI_sky130_fd_sc_hd__nor2_2
X_7655_ VGND VPWR _3075_ _3073_ _3074_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_141 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_7_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7586_ VGND VPWR _3012_ _3009_ _3011_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6606_ VPWR VGND VGND VPWR _3879_ _2054_ _2059_ _2060_ ZI_sky130_fd_sc_hd__nor3_2
XFILLER_0_62_526 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6537_ VGND VPWR VGND VPWR _1464_ _1341_ _1707_ _1672_ _1993_ _1386_ ZI_sky130_fd_sc_hd__a2111o_2
X_4798_ VPWR VGND VGND VPWR _0272_ _0204_ _3948_ _3900_ _4042_ _0273_ ZI_sky130_fd_sc_hd__a311o_2
XFILLER_0_70_570 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6468_ VGND VPWR VGND VPWR _1925_ _1924_ _1408_ _1350_ _1489_ _1424_ ZI_sky130_fd_sc_hd__a32o_2
X_6399_ _1523_ _1857_ _1289_ _1440_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5419_ VGND VPWR VGND VPWR _0888_ _0887_ _0684_ _0886_ ZI_sky130_fd_sc_hd__and3b_2
XFILLER_0_112_193 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8207_ VGND VPWR VGND VPWR _3548_ new_block[12] _3576_ _3573_ _1125_ _0119_ ZI_sky130_fd_sc_hd__o32a_2
X_8138_ VGND VPWR _3514_ _2626_ _3513_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8069_ VGND VPWR VGND VPWR _3152_ new_block[63] _3451_ _3449_ _2775_ _0106_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_85_607 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_69_147 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_38_523 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_38_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_61_581 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_110_119 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_68_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5770_ VGND VPWR _1234_ _0799_ _1188_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_534 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_90_109 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4721_ _3934_ _0197_ _3948_ _3946_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_4_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7440_ VGND VPWR VGND VPWR _2877_ _1193_ _2879_ _2878_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_71_312 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4652_ VGND VPWR _4189_ _4188_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_4_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7371_ VGND VPWR _2815_ _2810_ _2814_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4583_ VPWR VGND VPWR VGND _3945_ _4119_ _3893_ _4114_ _4120_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_52_570 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6322_ VGND VPWR VGND VPWR _1781_ _1775_ _1772_ _1780_ _1622_ ZI_sky130_fd_sc_hd__a211o_2
X_6253_ VPWR VGND VPWR VGND _1409_ _1408_ _1358_ _1378_ _1713_ ZI_sky130_fd_sc_hd__a22o_2
X_5204_ VGND VPWR _0674_ _0577_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6184_ VPWR VGND VPWR VGND _1379_ _1456_ _1394_ _1433_ _1645_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_35_3 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5135_ VGND VPWR VPWR VGND _0604_ _0603_ _0605_ _0551_ _3753_ ZI_sky130_fd_sc_hd__o211a_2
X_5066_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[106] sword_ctr_reg\[0\] _0536_
+ ZI_sky130_fd_sc_hd__or3_2
X_5968_ VPWR VGND VGND VPWR _1389_ _1430_ _1288_ ZI_sky130_fd_sc_hd__nor2_2
X_7707_ VGND VPWR _3123_ _4062_ _0376_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4919_ VGND VPWR VGND VPWR _4104_ new_block[100] _0392_ _0364_ _0362_ _0015_ ZI_sky130_fd_sc_hd__o32a_2
X_5899_ VGND VPWR _1361_ _1360_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7638_ VGND VPWR VGND VPWR _3059_ _0148_ _3060_ _3028_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_15_261 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7569_ VGND VPWR _2997_ _2799_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_101_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_58_607 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_58_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_81_654 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_34_570 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_108_296 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_80_175 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_79_28 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_21_220 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_80_197 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_21_242 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_95_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6940_ VGND VPWR VGND VPWR _2393_ _2162_ _2133_ _2105_ _2070_ ZI_sky130_fd_sc_hd__and4_2
X_6871_ VGND VPWR VGND VPWR _1911_ new_block[120] _2324_ _2321_ _2307_ _0035_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_88_253 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5822_ sword_ctr_reg\[1\] _1284_ sword_ctr_reg\[0\] new_block[16] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
X_5753_ VGND VPWR VGND VPWR _0748_ _0751_ _1214_ _1215_ _1217_ _1216_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_8_247 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4704_ VGND VPWR VPWR VGND _0178_ _0179_ _0176_ _0180_ ZI_sky130_fd_sc_hd__or3_2
X_8472_ VGND VPWR VPWR VGND clk _0074_ reset_n new_block[95] ZI_sky130_fd_sc_hd__dfrtp_2
X_5684_ VPWR VGND VPWR VGND _0964_ _0688_ _0963_ _0671_ _0702_ _1149_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_60_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7423_ VGND VPWR _2863_ _2860_ _2862_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_44_378 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4635_ VPWR VGND VGND VPWR _3993_ _4172_ _3933_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_71_164 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_8_53 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_25_592 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7354_ VGND VPWR _2800_ _2799_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4566_ VGND VPWR _4104_ _4103_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_12_253 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6305_ VGND VPWR _1765_ _1680_ _1764_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4497_ VGND VPWR VPWR VGND _3837_ _3885_ _3846_ _4035_ ZI_sky130_fd_sc_hd__or3_2
X_7285_ VGND VPWR _2733_ _0489_ _2732_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6236_ VGND VPWR VGND VPWR _1009_ new_block[113] _1696_ _1693_ _1675_ _0028_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_110_472 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6167_ VPWR VGND VPWR VGND _1625_ _1627_ _1626_ _1624_ _1628_ ZI_sky130_fd_sc_hd__or4_2
X_5118_ VPWR VGND _0586_ _0588_ _0587_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_6098_ VPWR VGND VPWR VGND _1554_ _1559_ _1556_ _1545_ _1560_ ZI_sky130_fd_sc_hd__or4_2
X_5049_ VPWR VGND VGND VPWR _0520_ _0516_ _0519_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_79_264 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_67_437 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_82_407 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_62_120 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_105_233 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_58_404 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_14_67 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_105_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_109_561 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_41_337 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4420_ VGND VPWR VPWR VGND _3955_ _3954_ _3958_ _3957_ _3956_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_111_225 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_111_203 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_1_445 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_22_584 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4351_ VPWR VGND VPWR VGND _3888_ _3889_ _3873_ _3875_ ZI_sky130_fd_sc_hd__or3b_2
X_7070_ _2126_ _2521_ _2186_ _2157_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_4282_ sword_ctr_reg\[1\] _3820_ sword_ctr_reg\[0\] new_block[7] VPWR VGND VPWR VGND
+ ZI_sky130_fd_sc_hd__and3_2
X_6021_ _1400_ _1483_ _1339_ _1408_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7972_ VPWR VGND VGND VPWR _3364_ _3358_ _3363_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_89_551 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_55_74 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6923_ VGND VPWR VGND VPWR _2172_ _2127_ _2174_ _2230_ _2376_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_36_109 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_64_407 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6854_ VGND VPWR _2308_ _4087_ _0447_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_278 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6785_ VPWR VGND _2070_ _2239_ _2175_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5805_ VGND VPWR VPWR VGND _1260_ _1267_ _1259_ _1268_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_57_470 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8524_ VGND VPWR VPWR VGND clk _0126_ reset_n new_block[19] ZI_sky130_fd_sc_hd__dfrtp_2
X_5736_ VPWR VGND VPWR VGND _0702_ _0929_ _0846_ _0546_ _1200_ ZI_sky130_fd_sc_hd__a22o_2
X_5667_ VPWR VGND _1133_ _1132_ _1058_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8455_ VGND VPWR VPWR VGND clk _0057_ reset_n new_block[78] ZI_sky130_fd_sc_hd__dfrtp_2
X_7406_ VGND VPWR _2847_ _1128_ _2846_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_44_197 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4618_ VPWR VGND VGND VPWR _4121_ _3976_ _4153_ _4141_ _4155_ _4154_ ZI_sky130_fd_sc_hd__o221a_2
XFILLER_0_60_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5598_ VGND VPWR _1065_ _0902_ _1064_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8386_ VGND VPWR VGND VPWR _3736_ _3734_ _0158_ _3738_ ZI_sky130_fd_sc_hd__a21o_2
X_7337_ VGND VPWR VGND VPWR _2784_ _2783_ _2782_ _2779_ ZI_sky130_fd_sc_hd__o21a_2
X_4549_ VGND VPWR _4087_ new_block[96] round_key[96] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7268_ VPWR VGND VPWR VGND _2228_ _2158_ _2302_ _2330_ _2716_ ZI_sky130_fd_sc_hd__a22o_2
X_6219_ VPWR VGND _1680_ round_key[30] new_block[30] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7199_ VPWR VGND _2229_ _2648_ _2159_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_23_337 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_50_134 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_51_646 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_106_564 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_31_370 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_25_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_98_392 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6570_ VGND VPWR VGND VPWR _2025_ _1427_ _1438_ _1782_ _2024_ ZI_sky130_fd_sc_hd__a211o_2
X_5521_ VGND VPWR _0989_ _0903_ _0988_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_164 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_27_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8240_ VPWR VGND _3606_ _0807_ _0808_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_26_197 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_42_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_112_501 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5452_ VGND VPWR _4103_ _4090_ _0921_ _0920_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
XFILLER_0_1_220 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_1_242 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5383_ _0698_ _0852_ _0582_ _0544_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8171_ VPWR VGND VGND VPWR _3544_ _3542_ _3543_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_112_545 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4403_ VGND VPWR _3941_ _3940_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4334_ VGND VPWR _3872_ _3871_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_112_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7122_ _2345_ _2572_ _2120_ _2188_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7053_ VGND VPWR VPWR VGND _2464_ _2503_ _2500_ _2504_ ZI_sky130_fd_sc_hd__or3_2
X_6004_ VGND VPWR _1466_ _1465_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4265_ VPWR VGND VGND VPWR _3802_ _3803_ _3796_ ZI_sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_19_Left_132 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7955_ VGND VPWR _3348_ _3344_ _3347_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_510 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7886_ VPWR VGND _3286_ block[110] round_key[110] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6906_ VPWR VGND VPWR VGND _2358_ _2194_ _2230_ _2327_ _2202_ _2359_ ZI_sky130_fd_sc_hd__a221o_2
X_6837_ VPWR VGND VPWR VGND _2177_ _2235_ _2114_ _2170_ _2291_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_77_598 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_18_632 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6768_ VGND VPWR _2222_ _2184_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8507_ VGND VPWR VPWR VGND clk _0109_ reset_n new_block[2] ZI_sky130_fd_sc_hd__dfrtp_2
X_5719_ VPWR VGND _1184_ _1071_ _0800_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_17_197 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_28_Left_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6699_ VPWR VGND VPWR VGND _2153_ _2125_ _2152_ ZI_sky130_fd_sc_hd__or2_2
X_8438_ VGND VPWR VPWR VGND clk _0040_ reset_n new_block[125] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_454 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8369_ VGND VPWR VGND VPWR _3640_ new_block[28] _3722_ _3720_ _2624_ _0135_ ZI_sky130_fd_sc_hd__o32a_2
XPHY_EDGE_ROW_37_Left_150 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_102_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_51_410 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_24_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_11_307 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_87_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_36_65 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_59_521 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4952_ VPWR VGND VPWR VGND _4189_ _3923_ _3845_ _3911_ _0425_ ZI_sky130_fd_sc_hd__a22o_2
X_7740_ VGND VPWR VGND VPWR _3153_ new_block[32] _3151_ _3147_ _4060_ _0075_ ZI_sky130_fd_sc_hd__o32a_2
X_4883_ VPWR VGND VPWR VGND _4042_ _3911_ _4002_ _4010_ _0357_ ZI_sky130_fd_sc_hd__a22o_2
X_7671_ VGND VPWR _3090_ _0148_ _0368_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_52_97 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6622_ VGND VPWR VGND VPWR sword_ctr_reg\[1\] sword_ctr_reg\[0\] new_block[89] _2076_
+ ZI_sky130_fd_sc_hd__nand3b_2
XFILLER_0_27_473 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_27_495 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_104_309 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6553_ VGND VPWR VGND VPWR _2009_ _2008_ _2007_ _2006_ ZI_sky130_fd_sc_hd__o21a_2
X_6484_ VPWR VGND VGND VPWR _1940_ _1939_ _1395_ _1368_ _1557_ _1941_ ZI_sky130_fd_sc_hd__a311o_2
X_5504_ VPWR VGND VPWR VGND _0971_ _0630_ _0778_ _0859_ _0712_ _0972_ ZI_sky130_fd_sc_hd__a221o_2
X_5435_ VPWR VGND _0904_ _0903_ _0801_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_112_331 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8223_ VPWR VGND _3591_ _0368_ _4069_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_112_353 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_65_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8154_ VGND VPWR VGND VPWR _3529_ _3528_ _3527_ _3524_ ZI_sky130_fd_sc_hd__o21a_2
X_5366_ VGND VPWR VGND VPWR _0835_ _0648_ _0654_ _0833_ _0834_ ZI_sky130_fd_sc_hd__a211o_2
X_5297_ VPWR VGND VGND VPWR _0632_ _0767_ _0687_ ZI_sky130_fd_sc_hd__nor2_2
X_8085_ VPWR VGND VGND VPWR _3466_ _3463_ _3465_ ZI_sky130_fd_sc_hd__nand2_2
X_4317_ VPWR VGND VGND VPWR _3854_ _3855_ _3849_ ZI_sky130_fd_sc_hd__nor2_2
X_7105_ VGND VPWR _2556_ new_block[99] round_key[99] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7036_ VGND VPWR _2488_ _2323_ _2487_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4248_ VGND VPWR VGND VPWR _0010_ _3785_ round[3] _3786_ _0000_ ZI_sky130_fd_sc_hd__a211o_2
X_7938_ VGND VPWR _3332_ _0371_ _0431_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7869_ VGND VPWR _3270_ _3047_ _3269_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_14_Right_14 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_108_637 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_92_365 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_21_605 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_33_498 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_20_137 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_103_386 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_23_Right_23 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_71_505 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_12_616 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5220_ VGND VPWR _0690_ _0668_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_11_159 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_41_Right_41 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5151_ VPWR VGND VGND VPWR _0621_ _0620_ _0579_ ZI_sky130_fd_sc_hd__nand2_2
X_5082_ VPWR VGND VGND VPWR new_block[76] sword_ctr_reg\[0\] _0552_ ZI_sky130_fd_sc_hd__or2b_2
XPHY_EDGE_ROW_50_Right_50 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5984_ VGND VPWR VPWR VGND _1318_ _1364_ _1352_ _1446_ ZI_sky130_fd_sc_hd__or3_2
X_7723_ VGND VPWR VPWR VGND _3136_ _3132_ _3138_ _3118_ _3137_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_19_237 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4935_ VGND VPWR VGND VPWR _0408_ _4181_ _3993_ _3999_ _3969_ _0407_ ZI_sky130_fd_sc_hd__o221ai_2
X_4866_ VGND VPWR VPWR VGND _0277_ _0339_ _0276_ _0340_ ZI_sky130_fd_sc_hd__or3_2
X_7654_ VGND VPWR _3074_ _4077_ _0143_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_153 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_7_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_27_281 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7585_ VGND VPWR _3011_ _2628_ _3010_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6605_ VGND VPWR VGND VPWR _3797_ _2055_ _2056_ _2057_ _2059_ _2058_ ZI_sky130_fd_sc_hd__o41ai_2
X_4797_ VGND VPWR VGND VPWR _4153_ _3854_ _0272_ _3961_ ZI_sky130_fd_sc_hd__a21oi_2
X_6536_ VGND VPWR VGND VPWR _1427_ _1619_ _1506_ _1553_ _1992_ _1991_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_105_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_42_262 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_70_582 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6467_ VPWR VGND VGND VPWR _1329_ _1363_ _1353_ _3755_ _1924_ ZI_sky130_fd_sc_hd__and4b_2
X_6398_ VPWR VGND VPWR VGND _1855_ _1376_ _1616_ _1340_ _1453_ _1856_ ZI_sky130_fd_sc_hd__a221o_2
X_5418_ VPWR VGND VGND VPWR _0567_ _0887_ _3880_ ZI_sky130_fd_sc_hd__nor2_2
X_8206_ VPWR VGND VPWR VGND _3575_ _3490_ _3574_ _3468_ _1898_ _3576_ ZI_sky130_fd_sc_hd__a221o_2
X_5349_ VPWR VGND VPWR VGND _4101_ _0524_ _0818_ _0816_ _0817_ _0819_ ZI_sky130_fd_sc_hd__a221o_2
X_8137_ VPWR VGND _3513_ _2695_ _1241_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8068_ VPWR VGND VPWR VGND _3149_ _3367_ _3450_ _3328_ _0902_ _3451_ ZI_sky130_fd_sc_hd__a221o_2
X_7019_ VGND VPWR VPWR VGND _2464_ _2470_ _2258_ _2471_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_38_557 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_93_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_110_109 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_61_593 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_84_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_84_630 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_29_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4720_ _4010_ _0196_ _3869_ _3910_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_56_365 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4651_ VPWR VGND VGND VPWR _3824_ _3844_ _3830_ _3863_ _4188_ ZI_sky130_fd_sc_hd__and4b_2
XFILLER_0_4_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_4_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7370_ VGND VPWR _2814_ _2811_ _2813_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4582_ VGND VPWR VGND VPWR _4115_ _4116_ _4119_ _3987_ ZI_sky130_fd_sc_hd__a21oi_2
X_6321_ VPWR VGND VPWR VGND _1776_ _1779_ _1777_ _1720_ _1780_ ZI_sky130_fd_sc_hd__or4_2
X_6252_ VPWR VGND VGND VPWR _1653_ _1712_ _1655_ ZI_sky130_fd_sc_hd__nor2_2
X_6183_ VPWR VGND VGND VPWR _1507_ _1644_ _1535_ ZI_sky130_fd_sc_hd__nor2_2
X_5203_ VGND VPWR VGND VPWR _0671_ _0669_ _0672_ _0673_ ZI_sky130_fd_sc_hd__a21o_2
X_5134_ VPWR VGND VGND VPWR _4097_ _0604_ new_block[108] ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_58_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5065_ VGND VPWR VPWR VGND sword_ctr_reg\[0\] _0535_ new_block[42] ZI_sky130_fd_sc_hd__and2b_2
XFILLER_0_28_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5967_ VGND VPWR VGND VPWR _1429_ _1427_ _1359_ _1341_ _1428_ _1424_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_109_209 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_75_641 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_35_505 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7706_ VGND VPWR VGND VPWR _2997_ new_block[93] _3122_ _3119_ _2686_ _0072_ ZI_sky130_fd_sc_hd__o32a_2
X_4918_ VPWR VGND VPWR VGND _4094_ _0391_ _0366_ _0390_ _0392_ ZI_sky130_fd_sc_hd__a22o_2
X_5898_ _1353_ _1360_ _1338_ _1319_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7637_ VGND VPWR _3059_ _3054_ _3058_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4849_ VPWR VGND VPWR VGND _3981_ _3934_ _4033_ _4002_ _3925_ _0323_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_62_346 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7568_ VPWR VGND VPWR VGND _2995_ _2960_ _2994_ _2984_ _0234_ _2996_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_99_81 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6519_ VPWR VGND VGND VPWR _1974_ _1483_ _1289_ _1332_ _1523_ _1975_ ZI_sky130_fd_sc_hd__a311o_2
XFILLER_0_15_273 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7499_ VGND VPWR _2933_ _1896_ _2932_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_97_221 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_78_490 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_108_231 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_65_162 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_81_666 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_34_560 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_110_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_80_187 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_21_254 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_21_276 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_95_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6870_ VPWR VGND VPWR VGND _1281_ _1909_ _2323_ _1959_ _2322_ _2324_ ZI_sky130_fd_sc_hd__a221o_2
X_5821_ VGND VPWR VGND VPWR _1283_ new_block[48] sword_ctr_reg\[1\] sword_ctr_reg\[0\]
+ ZI_sky130_fd_sc_hd__and3b_2
XFILLER_0_17_505 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5752_ VPWR VGND VPWR VGND _0846_ _0695_ _0602_ _0635_ _1216_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_57_641 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4703_ VGND VPWR VGND VPWR _3988_ _4021_ _0179_ _4181_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_60_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8471_ VGND VPWR VPWR VGND clk _0073_ reset_n new_block[94] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_72_655 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5683_ VPWR VGND VPWR VGND _1148_ _0667_ _0695_ ZI_sky130_fd_sc_hd__or2_2
X_7422_ VGND VPWR _2862_ _0805_ _2861_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4634_ VPWR VGND VGND VPWR _4110_ _4171_ _4153_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_12_210 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7353_ VGND VPWR _4099_ _3777_ _2799_ _3770_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
X_4565_ VGND VPWR _4099_ _3777_ _4103_ _4097_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
X_6304_ VPWR VGND _1764_ _1763_ _1762_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_69_73 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Right_4 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_12_265 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_100_92 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4496_ VPWR VGND VPWR VGND _4033_ _4019_ _3869_ _4009_ _4034_ ZI_sky130_fd_sc_hd__a22o_2
X_7284_ VGND VPWR _2732_ _2556_ _0523_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6235_ VPWR VGND VPWR VGND _1281_ _0524_ _1695_ _0816_ _1694_ _1696_ ZI_sky130_fd_sc_hd__a221o_2
X_6166_ VPWR VGND VGND VPWR _1462_ _1627_ _1460_ ZI_sky130_fd_sc_hd__nor2_2
X_6097_ VPWR VGND VPWR VGND _1558_ _1501_ _1531_ _1557_ _1523_ _1559_ ZI_sky130_fd_sc_hd__a221o_2
X_5117_ VPWR VGND VGND VPWR _3787_ _0567_ _0562_ _0587_ ZI_sky130_fd_sc_hd__nor3_2
X_5048_ VGND VPWR _0519_ _0517_ _0518_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6999_ VGND VPWR VGND VPWR _2279_ _2178_ _2450_ _2451_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_75_482 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_7_281 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_105_245 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_105_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_58_416 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_109_573 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_53_143 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_41_349 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4350_ VGND VPWR VGND VPWR _3882_ _3887_ _3877_ _3794_ _3865_ _3888_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_111_248 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4281_ VGND VPWR VPWR VGND sword_ctr_reg\[0\] _3819_ new_block[39] ZI_sky130_fd_sc_hd__and2b_2
X_6020_ VPWR VGND VGND VPWR _1466_ _1482_ _1385_ ZI_sky130_fd_sc_hd__nor2_2
X_7971_ VGND VPWR _3363_ _3360_ _3362_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6922_ VGND VPWR VGND VPWR _2375_ _2372_ _2136_ _2269_ _2374_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_49_449 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6853_ VPWR VGND VPWR VGND _2181_ _2306_ _2243_ _2153_ _2307_ ZI_sky130_fd_sc_hd__or4_2
X_5804_ VPWR VGND VPWR VGND _1261_ _1266_ _1264_ _0753_ _1267_ ZI_sky130_fd_sc_hd__or4_2
X_6784_ VGND VPWR VGND VPWR _2158_ _2236_ _2237_ _2238_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_71_96 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5735_ VGND VPWR VGND VPWR _1009_ new_block[109] _1199_ _1196_ _1181_ _0024_ ZI_sky130_fd_sc_hd__o32a_2
X_8523_ VGND VPWR VPWR VGND clk _0125_ reset_n new_block[18] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_346 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8454_ VGND VPWR VPWR VGND clk _0056_ reset_n new_block[77] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_95_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5666_ VPWR VGND _1132_ round_key[36] new_block[36] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7405_ VGND VPWR _2846_ _0912_ _2845_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4617_ VPWR VGND VGND VPWR _4154_ _3945_ _3845_ ZI_sky130_fd_sc_hd__nand2_2
X_5597_ VPWR VGND _1064_ round_key[59] new_block[59] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_102_226 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8385_ VPWR VGND VGND VPWR _3736_ _3737_ _3734_ ZI_sky130_fd_sc_hd__nor2_2
X_7336_ VGND VPWR VGND VPWR _2782_ _2779_ _2783_ _2642_ ZI_sky130_fd_sc_hd__a21oi_2
X_4548_ VGND VPWR VGND VPWR _4080_ _4071_ _4085_ _4086_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_40_393 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4479_ VGND VPWR VGND VPWR _4016_ _3969_ _4017_ _3962_ ZI_sky130_fd_sc_hd__a21oi_2
X_7267_ VGND VPWR VGND VPWR _2715_ _2073_ _2120_ _2507_ _2508_ ZI_sky130_fd_sc_hd__a211o_2
X_6218_ VGND VPWR _1679_ new_block[25] round_key[25] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7198_ VGND VPWR VGND VPWR _1911_ new_block[124] _2647_ _2644_ _2624_ _0039_ ZI_sky130_fd_sc_hd__o32a_2
X_6149_ VGND VPWR VGND VPWR _1490_ _1609_ _1447_ _1547_ _1610_ ZI_sky130_fd_sc_hd__o22a_2
XPHY_EDGE_ROW_79_Right_79 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_106_576 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Right_88 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_97_Right_97 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_58_246 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_27_611 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_39_493 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5520_ VPWR VGND _0988_ round_key[58] new_block[58] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_41_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_41_88 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_41_113 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5451_ VGND VPWR _0920_ round_key[105] new_block[105] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5382_ VPWR VGND _0600_ _0851_ _0650_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_8170_ VGND VPWR _3543_ _4078_ _3055_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4402_ VPWR VGND VPWR VGND _3901_ _3940_ _3830_ _3837_ ZI_sky130_fd_sc_hd__or3b_2
X_7121_ VPWR VGND _2189_ _2571_ _2157_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_4333_ VPWR VGND VPWR VGND _3863_ _3847_ _3824_ _3846_ _3871_ ZI_sky130_fd_sc_hd__or4_2
X_7052_ VPWR VGND VPWR VGND _2346_ _2502_ _2347_ _2257_ _2503_ ZI_sky130_fd_sc_hd__or4_2
X_4264_ VGND VPWR VGND VPWR _3797_ _3798_ _3799_ _3800_ _3802_ _3801_ ZI_sky130_fd_sc_hd__o41ai_2
X_6003_ VGND VPWR VPWR VGND _1352_ _1318_ _1382_ _1465_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_66_41 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_66_96 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7954_ VGND VPWR _3347_ _3345_ _3346_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6905_ _2192_ _2358_ _2186_ _2231_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7885_ VGND VPWR VPWR VGND _3283_ _3282_ _3285_ _3265_ _3284_ ZI_sky130_fd_sc_hd__o211a_2
X_6836_ VGND VPWR VGND VPWR _2290_ _2184_ _2193_ _2112_ ZI_sky130_fd_sc_hd__o21a_2
X_6767_ VGND VPWR VGND VPWR _2221_ _2214_ _2120_ _2217_ _2220_ ZI_sky130_fd_sc_hd__a211o_2
X_5718_ VGND VPWR _1183_ _1135_ _1182_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_154 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8506_ VGND VPWR VPWR VGND clk _0108_ reset_n new_block[1] ZI_sky130_fd_sc_hd__dfrtp_2
X_6698_ VGND VPWR VPWR VGND _2142_ _2151_ _2137_ _2152_ ZI_sky130_fd_sc_hd__or3_2
X_5649_ VPWR VGND VPWR VGND _1112_ _1114_ _1113_ _1111_ _1115_ ZI_sky130_fd_sc_hd__or4_2
X_8437_ VGND VPWR VPWR VGND clk _0039_ reset_n new_block[124] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_466 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8368_ VPWR VGND VPWR VGND _3521_ _4093_ _3721_ _0169_ _1885_ _3722_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_60_477 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7319_ VPWR VGND VPWR VGND _2260_ _2223_ _2208_ _2216_ _2766_ ZI_sky130_fd_sc_hd__a22o_2
X_8299_ VGND VPWR _3659_ _0907_ _1133_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_113 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_23_146 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_36_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4951_ VPWR VGND VGND VPWR _3906_ _3969_ _0424_ _3998_ _4023_ ZI_sky130_fd_sc_hd__o22ai_2
X_4882_ VGND VPWR VGND VPWR _3971_ _3976_ _0356_ _3882_ ZI_sky130_fd_sc_hd__a21oi_2
X_7670_ VGND VPWR _3089_ _3083_ _3088_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_430 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6621_ VGND VPWR VGND VPWR sword_ctr_reg\[0\] new_block[57] sword_ctr_reg\[1\] _2075_
+ ZI_sky130_fd_sc_hd__nand3b_2
X_6552_ VGND VPWR VGND VPWR _2007_ _2006_ _2008_ _1001_ ZI_sky130_fd_sc_hd__a21oi_2
X_6483_ _1354_ _1940_ _1395_ _1430_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_14_124 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5503_ VGND VPWR VGND VPWR _0633_ _0846_ _0970_ _0971_ ZI_sky130_fd_sc_hd__a21o_2
X_5434_ VPWR VGND _0903_ round_key[40] new_block[40] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_30_628 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8222_ VGND VPWR _3590_ _3586_ _3589_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_552 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_2_574 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8153_ VGND VPWR VGND VPWR _3527_ _3524_ _3528_ _3339_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_112_365 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7104_ VGND VPWR _2555_ _2549_ _2554_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5365_ _0592_ _0834_ _0698_ _0569_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_58_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8084_ VGND VPWR _3465_ _2972_ _3464_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5296_ VGND VPWR VGND VPWR _0766_ _0607_ _0765_ _0670_ ZI_sky130_fd_sc_hd__o21a_2
X_4316_ VGND VPWR _3854_ _3853_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7035_ VPWR VGND _2487_ _2421_ _2309_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4247_ VPWR VGND VGND VPWR _3785_ _3786_ round[3] ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_96_116 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7937_ VGND VPWR VGND VPWR _3331_ new_block[51] _3330_ _3327_ _1815_ _0094_ ZI_sky130_fd_sc_hd__o32a_2
X_7868_ VGND VPWR _3269_ _3043_ _3223_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6819_ VPWR VGND VGND VPWR _2054_ _2273_ _3776_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_9_162 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7799_ VPWR VGND VGND VPWR _3207_ _3201_ _3206_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_107_137 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_21_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_60_274 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_68_330 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Left_114 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_56_514 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_43_208 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_43_219 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_12_628 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_51_241 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_106_181 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5150_ VGND VPWR _0620_ _0598_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5081_ VGND VPWR VGND VPWR _0538_ _0547_ _0548_ _0549_ _0550_ _0551_ ZI_sky130_fd_sc_hd__o41a_2
XFILLER_0_47_43 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_47_98 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_79_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5983_ VPWR VGND VGND VPWR _1445_ _1444_ _1368_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_78_149 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Left_169 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4934_ VGND VPWR VGND VPWR _3941_ _3954_ _3992_ _3930_ _3948_ _0407_ ZI_sky130_fd_sc_hd__o32a_2
X_7722_ VPWR VGND VGND VPWR _3137_ _3132_ _3136_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_7_600 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_74_322 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4865_ VGND VPWR VGND VPWR _0338_ _0337_ _0339_ _0336_ _0335_ ZI_sky130_fd_sc_hd__nand4_2
X_7653_ VGND VPWR _3073_ _0298_ _0380_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_121 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7584_ VGND VPWR _3010_ _2011_ _2490_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6604_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[124] sword_ctr_reg\[0\] _2058_
+ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_74_377 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4796_ VGND VPWR _0270_ _3949_ _0271_ _0268_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
X_6535_ VPWR VGND VPWR VGND _1361_ _1452_ _1345_ _1499_ _1991_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_70_550 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_15_499 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6466_ VPWR VGND VPWR VGND _1350_ _1426_ _1359_ _1397_ _1923_ ZI_sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_65_Left_178 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8205_ VGND VPWR _3575_ _3458_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6397_ VPWR VGND VGND VPWR _1552_ _1855_ _1385_ ZI_sky130_fd_sc_hd__nor2_2
X_5417_ VPWR VGND VGND VPWR _0562_ _0886_ _3880_ ZI_sky130_fd_sc_hd__nor2_2
X_5348_ VPWR VGND _0818_ new_block[104] round_key[104] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8136_ VGND VPWR _3512_ _2776_ _3511_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8067_ VPWR VGND _3450_ block[63] round_key[63] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7018_ VGND VPWR VGND VPWR _2470_ _2222_ _2194_ _2467_ _2469_ ZI_sky130_fd_sc_hd__a211o_2
X_5279_ VGND VPWR VGND VPWR _0749_ _0569_ _0596_ _0684_ _0705_ ZI_sky130_fd_sc_hd__and4_2
XPHY_EDGE_ROW_74_Left_187 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_77_182 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_65_322 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_38_569 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_93_653 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_92_141 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_53_517 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_65_388 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_18_282 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_33_263 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_83_Left_196 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_61_561 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_103_162 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_103_184 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_108_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4650_ VPWR VGND VGND VPWR _3965_ _4187_ _3898_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_4_625 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6320_ VGND VPWR VGND VPWR _1779_ _1397_ _1778_ _1464_ ZI_sky130_fd_sc_hd__o21a_2
X_4581_ VGND VPWR VGND VPWR _4118_ _3955_ _4115_ _3954_ _4114_ _4117_ ZI_sky130_fd_sc_hd__o221ai_2
XFILLER_0_71_369 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_52_583 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6251_ VPWR VGND VPWR VGND _1708_ _1710_ _1709_ _1707_ _1711_ ZI_sky130_fd_sc_hd__or4_2
X_6182_ VPWR VGND VGND VPWR _1628_ _1634_ _1642_ _1643_ ZI_sky130_fd_sc_hd__nor3_2
X_5202_ VGND VPWR VGND VPWR _0672_ _0600_ _0557_ _0582_ _0620_ ZI_sky130_fd_sc_hd__and4_2
X_5133_ VPWR VGND VPWR VGND _0552_ _3764_ _0603_ _0553_ _0554_ ZI_sky130_fd_sc_hd__a211oi_2
XFILLER_0_74_41 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5064_ sword_ctr_reg\[1\] _0534_ sword_ctr_reg\[0\] new_block[10] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_79_403 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_74_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_94_417 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_66_108 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5966_ _1295_ _1428_ _1400_ _1369_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5897_ VGND VPWR _1359_ _1358_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7705_ VGND VPWR VGND VPWR _3122_ _3120_ _4094_ _3121_ _2797_ ZI_sky130_fd_sc_hd__a211o_2
X_4917_ VPWR VGND _0391_ block[68] round_key[68] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_74_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7636_ VGND VPWR _3058_ _3056_ _3057_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4848_ VPWR VGND VPWR VGND _0265_ _3900_ _4042_ _4012_ _4019_ _0322_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_28_580 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_90_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4779_ VPWR VGND VGND VPWR _4021_ _0254_ _3987_ ZI_sky130_fd_sc_hd__nor2_2
X_7567_ VGND VPWR _2995_ _2796_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6518_ _1354_ _1974_ _1289_ _1437_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_99_93 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7498_ VGND VPWR _2932_ _1833_ _2003_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6449_ VPWR VGND _1907_ block[20] round_key[20] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_100_132 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8119_ VPWR VGND VGND VPWR _3496_ _3497_ _3495_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_97_277 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_38_344 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_108_221 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_91_Left_204 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_1_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_88_222 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5820_ VGND VPWR VGND VPWR _1009_ new_block[111] _1282_ _1278_ _1268_ _0026_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_48_119 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5751_ VPWR VGND VPWR VGND _0580_ _0571_ _0613_ _0607_ _1215_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_84_450 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_60_21 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_56_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_29_388 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4702_ VGND VPWR VGND VPWR _0178_ _3924_ _0177_ _4010_ _3911_ _3894_ ZI_sky130_fd_sc_hd__a32o_2
X_8470_ VGND VPWR VPWR VGND clk _0072_ reset_n new_block[93] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_72_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5682_ VGND VPWR VGND VPWR _1009_ new_block[108] _1147_ _1144_ _1125_ _0023_ ZI_sky130_fd_sc_hd__o32a_2
X_7421_ VPWR VGND _2861_ _0902_ _0811_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_71_122 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_60_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_25_561 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4633_ VPWR VGND VPWR VGND _3900_ _4033_ _3923_ _3925_ _4170_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_72_667 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_102_408 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7352_ VPWR VGND VPWR VGND _2797_ _2786_ _2795_ _2703_ _0147_ _2798_ ZI_sky130_fd_sc_hd__a221o_2
X_4564_ VGND VPWR VGND VPWR _4101_ _4094_ _4095_ _4096_ _4102_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_12_222 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7283_ VGND VPWR VGND VPWR _2731_ _3756_ _2730_ _2708_ ZI_sky130_fd_sc_hd__o21a_2
X_6303_ VPWR VGND _1763_ round_key[26] new_block[26] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6234_ VPWR VGND _1695_ new_block[113] round_key[113] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4495_ _3891_ _4033_ _3831_ _3901_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6165_ VPWR VGND _1474_ _1626_ _1396_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_40_3 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_85_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6096_ VPWR VGND _1491_ _1558_ _1409_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5116_ VGND VPWR VGND VPWR _0586_ _0556_ _0555_ _0551_ _3753_ ZI_sky130_fd_sc_hd__and4_2
X_5047_ VPWR VGND _0518_ _0383_ _0150_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6998_ _2173_ _2450_ _2188_ _2368_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5949_ VGND VPWR VGND VPWR _1411_ _1403_ _1390_ _1406_ _1410_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_62_100 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_7_271 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7619_ VGND VPWR VGND VPWR _2997_ new_block[86] _3042_ _3040_ _1996_ _0065_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_63_667 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_90_497 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_98_542 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_105_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_38_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_109_541 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_38_174 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_81_431 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_66_494 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_54_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_54_634 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_109_585 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4280_ VPWR VGND VGND VPWR new_block[71] sword_ctr_reg\[0\] _3818_ ZI_sky130_fd_sc_hd__or2b_2
X_7970_ VGND VPWR _3362_ _3111_ _3361_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_87 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6921_ VPWR VGND VPWR VGND _2190_ _2373_ _2115_ _2168_ _2374_ ZI_sky130_fd_sc_hd__a22o_2
X_6852_ VPWR VGND VPWR VGND _2277_ _2305_ _2293_ _2251_ _2306_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_76_203 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5803_ VGND VPWR VGND VPWR _1266_ _0727_ _0726_ _1164_ _1265_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_71_53 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8522_ VGND VPWR VPWR VGND clk _0124_ reset_n new_block[17] ZI_sky130_fd_sc_hd__dfrtp_2
X_6783_ VGND VPWR VGND VPWR _2237_ _2199_ _2161_ _2070_ _2182_ ZI_sky130_fd_sc_hd__and4_2
X_5734_ VPWR VGND VPWR VGND _4101_ _0524_ _1198_ _0816_ _1197_ _1199_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_29_185 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5665_ VGND VPWR _1131_ _0795_ _0909_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_44_155 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_44_166 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8453_ VGND VPWR VPWR VGND clk _0055_ reset_n new_block[76] ZI_sky130_fd_sc_hd__dfrtp_2
X_7404_ VPWR VGND _2845_ _1068_ _0992_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8384_ VGND VPWR _3736_ _2953_ _3735_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_60_637 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4616_ VPWR VGND VGND VPWR _4153_ _3869_ _3959_ ZI_sky130_fd_sc_hd__nand2_2
X_5596_ VPWR VGND _1063_ _0993_ _0810_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7335_ VGND VPWR _2782_ _2694_ _2781_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_111_Right_111 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_111_81 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_4_296 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_102_238 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4547_ VGND VPWR _4085_ _4084_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4478_ VPWR VGND VGND VPWR _4016_ _3815_ _3959_ ZI_sky130_fd_sc_hd__nand2_2
X_7266_ VGND VPWR VPWR VGND _2711_ _2713_ _2582_ _2714_ ZI_sky130_fd_sc_hd__or3_2
X_7197_ VPWR VGND VPWR VGND _4100_ _1909_ _2646_ _1959_ _2645_ _2647_ ZI_sky130_fd_sc_hd__a221o_2
X_6217_ VGND VPWR _1678_ _1564_ _1677_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6148_ VGND VPWR _1609_ _1608_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6079_ VPWR VGND VPWR VGND _1526_ _1540_ _1533_ _1520_ _1541_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_67_225 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_36_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_23_306 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_35_133 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_35_144 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_106_533 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_35_177 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_90_261 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_42_604 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_54_442 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5450_ VPWR VGND VPWR VGND _0919_ round_key[41] block[41] ZI_sky130_fd_sc_hd__or2_2
XFILLER_0_41_125 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_41_136 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4401_ VGND VPWR VGND VPWR _3749_ _3751_ _3793_ _3802_ _3910_ _3939_ ZI_sky130_fd_sc_hd__o41a_2
XFILLER_0_41_169 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5381_ VPWR VGND VPWR VGND _0785_ _0546_ _0705_ _0589_ _0850_ ZI_sky130_fd_sc_hd__a22o_2
X_7120_ VGND VPWR VGND VPWR _2360_ _2127_ _2567_ _2568_ _2570_ _2569_ ZI_sky130_fd_sc_hd__a2111o_2
X_4332_ VPWR VGND VGND VPWR _3870_ _3804_ _3869_ ZI_sky130_fd_sc_hd__nand2_2
X_4263_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[97] sword_ctr_reg\[0\] _3801_
+ ZI_sky130_fd_sc_hd__or3_2
X_7051_ VGND VPWR VGND VPWR _2435_ _2166_ _2501_ _2502_ ZI_sky130_fd_sc_hd__a21o_2
X_6002_ VPWR VGND VGND VPWR _1455_ _1464_ _1307_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_66_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7953_ VGND VPWR _3346_ _0239_ _0385_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_309 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_82_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_49_203 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6904_ VPWR VGND VPWR VGND _2353_ _2356_ _2354_ _2352_ _2357_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_77_501 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_49_225 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_49_258 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7884_ VPWR VGND VGND VPWR _3284_ _3282_ _3283_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_106_81 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_82_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_92_526 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6835_ VGND VPWR VGND VPWR _2289_ _2112_ _2281_ _2101_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_18_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_45_420 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6766_ VPWR VGND VPWR VGND _2219_ _2218_ _2214_ _2155_ _2220_ ZI_sky130_fd_sc_hd__a22o_2
X_5717_ VGND VPWR _1182_ _0811_ _1065_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_388 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8505_ VGND VPWR VPWR VGND clk _0107_ reset_n new_block[0] ZI_sky130_fd_sc_hd__dfrtp_2
X_6697_ VPWR VGND VPWR VGND _2150_ _2149_ _2073_ _2144_ _2151_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_32_136 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8436_ VGND VPWR VPWR VGND clk _0038_ reset_n new_block[123] ZI_sky130_fd_sc_hd__dfrtp_2
X_5648_ VPWR VGND VPWR VGND _0627_ _0731_ _0606_ _0729_ _1114_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_20_309 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8367_ VPWR VGND _3721_ block[28] round_key[28] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_60_489 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5579_ VGND VPWR VGND VPWR _1046_ _0825_ _0648_ _0616_ ZI_sky130_fd_sc_hd__o21a_2
X_8298_ VGND VPWR VGND VPWR _3640_ new_block[21] _3658_ _3656_ _1943_ _0128_ ZI_sky130_fd_sc_hd__o32a_2
X_7318_ VGND VPWR VGND VPWR _2765_ _2246_ _2107_ _2389_ _2423_ ZI_sky130_fd_sc_hd__a211o_2
X_7249_ VGND VPWR _2698_ _2693_ _2697_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_125 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_68_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_24_615 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_78_309 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_59_534 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4950_ VGND VPWR VGND VPWR _0418_ _4008_ _0420_ _0343_ _0423_ _0422_ ZI_sky130_fd_sc_hd__a2111o_2
X_4881_ VGND VPWR VGND VPWR _3969_ _4021_ _0355_ _3962_ ZI_sky130_fd_sc_hd__a21oi_2
X_6620_ VGND VPWR VGND VPWR new_block[25] sword_ctr_reg\[0\] _2074_ sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__nand3_2
XFILLER_0_74_559 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6551_ VGND VPWR _2007_ _1892_ _1945_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5502_ VGND VPWR VGND VPWR _0970_ _0569_ _0592_ _0583_ _0532_ ZI_sky130_fd_sc_hd__and4_2
X_6482_ VGND VPWR VGND VPWR _1938_ _1447_ _1939_ _1404_ ZI_sky130_fd_sc_hd__a21oi_2
X_5433_ VPWR VGND _0902_ round_key[63] new_block[63] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8221_ VGND VPWR _3589_ _0485_ _3588_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5364_ VGND VPWR VGND VPWR _0833_ _0569_ _0545_ _0698_ _0532_ ZI_sky130_fd_sc_hd__and4_2
X_8152_ VGND VPWR _3527_ _2637_ _3526_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7103_ VGND VPWR _2554_ _2551_ _2553_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4315_ VGND VPWR VPWR VGND _3794_ _3852_ _3851_ _3853_ ZI_sky130_fd_sc_hd__or3_2
X_5295_ _0577_ _0765_ _0531_ _0579_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8083_ VGND VPWR _3464_ _2308_ _2630_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7034_ VGND VPWR _2486_ _0818_ _1241_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4246_ VGND VPWR VGND VPWR _3748_ keylen _3785_ _0009_ _3784_ ZI_sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_93_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_96_106 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7936_ VGND VPWR _3331_ _3152_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7867_ VGND VPWR VGND VPWR _3240_ new_block[44] _3268_ _3266_ _1125_ _0087_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_9_130 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6818_ VPWR VGND VPWR VGND _2195_ _2264_ _2141_ _2167_ _2272_ ZI_sky130_fd_sc_hd__a22o_2
X_7798_ VGND VPWR _3206_ _3203_ _3205_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_107_149 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6749_ VGND VPWR _2203_ _2162_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_45_294 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8419_ VGND VPWR VPWR VGND clk _0021_ reset_n new_block[106] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_21_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_103_333 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_13_191 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_83_389 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_71_518 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_98_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_106_193 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_11_106 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_102_Left_215 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5080_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[109] sword_ctr_reg\[0\] _0550_
+ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_79_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5982_ VGND VPWR _1444_ _1441_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4933_ VPWR VGND VPWR VGND _0178_ _0405_ _0404_ _3855_ _0406_ ZI_sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_111_Left_224 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7721_ VGND VPWR _3136_ _3133_ _3135_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_515 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_7_612 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4864_ VGND VPWR VGND VPWR _3872_ _3921_ _3974_ _4036_ _0338_ ZI_sky130_fd_sc_hd__o22a_2
X_7652_ VGND VPWR VGND VPWR _2997_ new_block[89] _3072_ _3070_ _2408_ _0068_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_6_133 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_27_272 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7583_ VPWR VGND _3009_ _2738_ _2646_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4795_ VPWR VGND VGND VPWR _4141_ _3816_ _3998_ _3870_ _0270_ _0269_ ZI_sky130_fd_sc_hd__o221a_2
XFILLER_0_105_609 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6603_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] _2057_ new_block[92] ZI_sky130_fd_sc_hd__and2b_2
X_6534_ VGND VPWR VGND VPWR _1606_ _1515_ _1987_ _1988_ _1990_ _1989_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_55_592 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6465_ VPWR VGND VPWR VGND _1921_ _1633_ _1922_ _1439_ _1638_ ZI_sky130_fd_sc_hd__or4b_2
X_5416_ VGND VPWR VGND VPWR _0885_ _0689_ _0669_ _0627_ ZI_sky130_fd_sc_hd__o21a_2
X_8204_ VPWR VGND _3574_ block[76] round_key[76] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_112_141 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6396_ VGND VPWR VGND VPWR _1854_ _1431_ _1379_ _1515_ _1602_ _1395_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_100_303 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5347_ VPWR VGND _0817_ block[40] round_key[40] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8135_ VPWR VGND _3511_ _2625_ _2310_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8066_ VGND VPWR VPWR VGND _3446_ _3445_ _3449_ _3448_ _3447_ ZI_sky130_fd_sc_hd__o211a_2
X_5278_ VGND VPWR _0748_ _0713_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7017_ VGND VPWR VGND VPWR _2468_ _2343_ _2229_ _2214_ _2469_ ZI_sky130_fd_sc_hd__a31o_2
X_4229_ VPWR VGND VGND VPWR dec_ctrl_reg\[3\] _3772_ dec_ctrl_reg\[2\] ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_69_106 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_78_640 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_69_139 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7919_ VGND VPWR _3315_ _0232_ _0299_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_161 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_46_570 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_80_359 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_21_404 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_61_551 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_103_152 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_103_196 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_88_459 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_88_448 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_75_109 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_33_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4580_ VGND VPWR VGND VPWR _4023_ _4116_ _4114_ _4117_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_4_637 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_24_253 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_109_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6250_ VGND VPWR VGND VPWR _1440_ _1527_ _1539_ _1536_ _1710_ _1544_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_110_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6181_ VGND VPWR VPWR VGND _1638_ _1641_ _1423_ _1642_ ZI_sky130_fd_sc_hd__or3_2
X_5201_ VGND VPWR _0671_ _0670_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_110_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5132_ VGND VPWR _0602_ _0601_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5063_ VGND VPWR VGND VPWR _0533_ sword_ctr_reg\[0\] new_block[74] sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__and3b_2
XFILLER_0_74_97 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_94_407 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5965_ VGND VPWR _1427_ _1426_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_90_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5896_ VPWR VGND VGND VPWR _1357_ _1358_ _1295_ ZI_sky130_fd_sc_hd__nor2_2
X_4916_ VGND VPWR _0390_ _0372_ _0389_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7704_ VPWR VGND VGND VPWR _4062_ _3121_ _4090_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_35_518 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_47_389 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4847_ VGND VPWR VPWR VGND _0175_ _0180_ _3980_ _0321_ ZI_sky130_fd_sc_hd__or3_2
X_7635_ VGND VPWR _3057_ _4078_ _0153_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_475 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_90_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_74_197 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_7_497 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7566_ VPWR VGND _2994_ block[114] round_key[114] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4778_ VPWR VGND VPWR VGND _3920_ _4143_ _4033_ _4003_ _0253_ ZI_sky130_fd_sc_hd__a22o_2
X_6517_ VGND VPWR VPWR VGND _1964_ _1972_ _1648_ _1973_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_43_573 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7497_ VGND VPWR _2931_ _2927_ _2930_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6448_ VGND VPWR VGND VPWR _1906_ _1905_ _1904_ _1893_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_100_111 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6379_ VGND VPWR VGND VPWR _1837_ _1827_ _1838_ _1001_ ZI_sky130_fd_sc_hd__a21oi_2
X_8118_ VGND VPWR _3496_ _2417_ _3026_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8049_ VPWR VGND VGND VPWR _3433_ round_key[62] block[62] ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_26_529 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_93_462 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_1_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_88_234 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_88_212 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_69_470 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5750_ VPWR VGND VPWR VGND _0729_ _0635_ _0613_ _0627_ _1214_ ZI_sky130_fd_sc_hd__a22o_2
X_5681_ VPWR VGND VPWR VGND _4101_ _0524_ _1146_ _0816_ _1145_ _1147_ ZI_sky130_fd_sc_hd__a221o_2
X_4701_ VPWR VGND VGND VPWR _3878_ _0177_ _3794_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_84_462 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_72_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_57_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_56_164 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7420_ VGND VPWR _2860_ _0800_ _1139_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_44_348 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4632_ VGND VPWR VGND VPWR _4042_ _4168_ _3988_ _3887_ _4169_ ZI_sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_56_197 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_60_99 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7351_ VGND VPWR _2797_ _2796_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4563_ VGND VPWR _4101_ _4100_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_12_234 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7282_ VPWR VGND VPWR VGND _2718_ _2729_ _2726_ _2714_ _2730_ ZI_sky130_fd_sc_hd__or4_2
X_6302_ VPWR VGND _1762_ round_key[31] new_block[31] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4494_ VPWR VGND VPWR VGND _3903_ _4031_ _3911_ _4030_ _4032_ ZI_sky130_fd_sc_hd__a22o_2
X_6233_ VPWR VGND _1694_ block[17] round_key[17] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_12_278 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6164_ VPWR VGND VGND VPWR _1462_ _1625_ _1370_ ZI_sky130_fd_sc_hd__nor2_2
X_6095_ VGND VPWR _1557_ _1499_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_85_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5115_ VGND VPWR VGND VPWR _0584_ _0546_ _0585_ _0571_ ZI_sky130_fd_sc_hd__a21bo_2
XFILLER_0_33_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_109_81 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5046_ VGND VPWR _0517_ _4069_ _0431_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_96 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6997_ VGND VPWR VGND VPWR _2449_ _2282_ _2256_ _2447_ _2448_ ZI_sky130_fd_sc_hd__a211o_2
X_5948_ _1408_ _1410_ _1400_ _1409_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_94_237 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5879_ VGND VPWR _1341_ _1340_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7618_ VPWR VGND VPWR VGND _2995_ _3041_ _2857_ _2984_ _4073_ _3042_ ZI_sky130_fd_sc_hd__a221o_2
X_7549_ VGND VPWR _2978_ _2550_ _2552_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_475 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_14_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_105_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_38_164 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_39_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_38_186 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_53_123 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_109_553 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_93_281 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_66_484 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_109_597 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_54_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6920_ VGND VPWR _2373_ _2176_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6851_ VPWR VGND VPWR VGND _2296_ _2304_ _2298_ _2295_ _2305_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_89_587 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_9_526 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5802_ VPWR VGND VPWR VGND _0870_ _0846_ _0975_ _0616_ _0658_ _1265_ ZI_sky130_fd_sc_hd__a221o_2
X_8521_ VGND VPWR VPWR VGND clk _0123_ reset_n new_block[16] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_602 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6782_ VGND VPWR _2236_ _2235_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5733_ VPWR VGND _1198_ new_block[109] round_key[109] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_45_635 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_84_281 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_72_421 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5664_ VPWR VGND _1130_ _1129_ _1127_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_44_134 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8452_ VGND VPWR VPWR VGND clk _0054_ reset_n new_block[75] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_242 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5595_ VGND VPWR _1062_ _0998_ _1061_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8383_ VPWR VGND _3735_ _3202_ _1898_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4615_ VPWR VGND VPWR VGND _4151_ _4047_ _3931_ _3910_ _4152_ ZI_sky130_fd_sc_hd__a22o_2
X_7403_ VGND VPWR VGND VPWR _2800_ new_block[68] _2844_ _2842_ _0362_ _0047_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_4_253 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7334_ VGND VPWR _2781_ _2048_ _2780_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4546_ VPWR VGND VPWR VGND _4084_ _4082_ _4083_ ZI_sky130_fd_sc_hd__or2_2
XFILLER_0_111_93 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4477_ VPWR VGND VGND VPWR _3987_ _4015_ _3854_ ZI_sky130_fd_sc_hd__nor2_2
X_7265_ VGND VPWR VGND VPWR _2713_ _2360_ _2219_ _2605_ _2712_ ZI_sky130_fd_sc_hd__a211o_2
X_7196_ VPWR VGND _2646_ new_block[124] round_key[124] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6216_ VPWR VGND _1677_ _1676_ _1569_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6147_ VGND VPWR VPWR VGND _1363_ _1364_ _1313_ _1608_ ZI_sky130_fd_sc_hd__or3_2
X_6078_ VGND VPWR VGND VPWR _1536_ _1534_ _1539_ _1540_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_99_329 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5029_ VPWR VGND VPWR VGND _3947_ _3986_ _0499_ _3897_ _0500_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_95_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_36_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_8_581 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_106_545 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_90_273 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_106_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_58_215 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_26_101 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_42_616 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4400_ VPWR VGND VGND VPWR _3905_ _3938_ _3877_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_1_234 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5380_ VGND VPWR VGND VPWR _0849_ _0667_ _0662_ _0673_ _0641_ ZI_sky130_fd_sc_hd__a211o_2
X_4331_ VGND VPWR _3869_ _3868_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4262_ VGND VPWR VGND VPWR _3800_ sword_ctr_reg\[0\] new_block[65] sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__and3b_2
X_7050_ VGND VPWR VGND VPWR _2501_ _2256_ _2222_ _2196_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_5_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6001_ VGND VPWR VGND VPWR _1460_ _1412_ _1463_ _1462_ ZI_sky130_fd_sc_hd__a21oi_2
X_7952_ VGND VPWR _3345_ _4073_ _0309_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_215 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6903_ VGND VPWR VGND VPWR _2356_ _2300_ _2223_ _2355_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_82_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7883_ VGND VPWR _3283_ _2646_ _2739_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6834_ VPWR VGND VPWR VGND _2106_ _2157_ _2101_ _2201_ _2288_ ZI_sky130_fd_sc_hd__a22o_2
X_6765_ VGND VPWR _2219_ _2188_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_18_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8504_ VGND VPWR VPWR VGND clk _0106_ reset_n new_block[63] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_432 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5716_ VPWR VGND VPWR VGND _1157_ _1180_ _1160_ _1156_ _1181_ ZI_sky130_fd_sc_hd__or4_2
X_8435_ VGND VPWR VPWR VGND clk _0037_ reset_n new_block[122] ZI_sky130_fd_sc_hd__dfrtp_2
X_6696_ VGND VPWR _2150_ _2101_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5647_ VPWR VGND VGND VPWR _0948_ _1113_ _0640_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_60_435 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8366_ VGND VPWR VPWR VGND _3718_ _1897_ _3720_ _0366_ _3719_ ZI_sky130_fd_sc_hd__o211a_2
X_5578_ VGND VPWR VGND VPWR _1041_ _0923_ _1044_ _1045_ ZI_sky130_fd_sc_hd__a21o_2
X_8297_ VPWR VGND VPWR VGND _3575_ _3603_ _3657_ _3583_ _1569_ _3658_ ZI_sky130_fd_sc_hd__a221o_2
X_7317_ VPWR VGND VPWR VGND _2168_ _2282_ _2256_ _2178_ _2764_ ZI_sky130_fd_sc_hd__a22o_2
X_4529_ VPWR VGND _4067_ round_key[70] new_block[70] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7248_ VGND VPWR _2697_ _2694_ _2696_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7179_ VGND VPWR _2629_ _2627_ _2628_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_137 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_68_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_11_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_24_627 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_36_487 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_102_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_102_581 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_59_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_59_546 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4880_ VGND VPWR VGND VPWR _4021_ _4115_ _0354_ _4110_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_39_281 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6550_ VGND VPWR _2006_ _1999_ _2005_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5501_ VGND VPWR VGND VPWR _0969_ _0888_ _0671_ _0965_ _0968_ ZI_sky130_fd_sc_hd__a211o_2
X_6481_ VPWR VGND VGND VPWR _1938_ _1313_ _1414_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_14_148 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5432_ VGND VPWR _0901_ _0805_ _0900_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8220_ VGND VPWR _3588_ _0382_ _3587_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8151_ VGND VPWR _3526_ _3033_ _3525_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5363_ VPWR VGND VPWR VGND _0824_ _0831_ _0830_ _0821_ _0832_ ZI_sky130_fd_sc_hd__or4_2
X_7102_ VPWR VGND _2553_ _2552_ _2490_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4314_ VPWR VGND VPWR VGND _3852_ _3832_ _3802_ ZI_sky130_fd_sc_hd__or2_2
X_8082_ VPWR VGND _3463_ _2546_ _2409_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5294_ VPWR VGND VPWR VGND _0656_ _0763_ _0664_ _0690_ _0764_ ZI_sky130_fd_sc_hd__a22o_2
X_7033_ VPWR VGND _2485_ _2484_ _0489_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4245_ VPWR VGND VPWR VGND _3785_ round[2] _3782_ ZI_sky130_fd_sc_hd__or2_2
X_7935_ VPWR VGND VPWR VGND _3309_ _3257_ _3329_ _3328_ _1068_ _3330_ ZI_sky130_fd_sc_hd__a221o_2
X_7866_ VPWR VGND VPWR VGND _3219_ _3257_ _3267_ _3237_ _1188_ _3268_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_65_505 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6817_ VPWR VGND _2134_ _2271_ _2201_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_92_357 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7797_ VPWR VGND _3205_ _3204_ _2912_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6748_ VGND VPWR _2202_ _2201_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6679_ VPWR VGND VGND VPWR _3787_ _2133_ _2059_ _2054_ ZI_sky130_fd_sc_hd__nor3b_2
XFILLER_0_60_221 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8418_ VGND VPWR VPWR VGND clk _0020_ reset_n new_block[105] ZI_sky130_fd_sc_hd__dfrtp_2
X_8349_ VPWR VGND VPWR VGND _3521_ _3603_ _3704_ _0169_ _1763_ _3705_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_96_641 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_68_365 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_56_527 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_49_590 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_106_150 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_51_298 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_10_Right_10 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5981_ VGND VPWR _1443_ _1442_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_87_630 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_47_505 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7720_ VGND VPWR _3135_ _0437_ _3134_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4932_ VGND VPWR VGND VPWR _0405_ _4041_ _3997_ _4189_ _4003_ _3795_ ZI_sky130_fd_sc_hd__a32o_2
X_7651_ VPWR VGND VPWR VGND _2995_ _2960_ _3071_ _2984_ _0143_ _3072_ ZI_sky130_fd_sc_hd__a221o_2
X_4863_ VGND VPWR VPWR VGND _3939_ _3992_ _3930_ _0337_ ZI_sky130_fd_sc_hd__or3_2
X_6602_ sword_ctr_reg\[1\] _2056_ sword_ctr_reg\[0\] new_block[28] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
X_7582_ VGND VPWR _3008_ _2485_ _2638_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4794_ VGND VPWR VGND VPWR _3998_ _0182_ _4052_ _4131_ _0269_ ZI_sky130_fd_sc_hd__o22a_2
X_6533_ VPWR VGND VPWR VGND _1470_ _1529_ _1351_ _1531_ _1989_ ZI_sky130_fd_sc_hd__a22o_2
X_6464_ VPWR VGND VPWR VGND _1811_ _1603_ _1525_ _1422_ _1921_ ZI_sky130_fd_sc_hd__or4_2
X_5415_ VPWR VGND VPWR VGND _0883_ _0709_ _0701_ _0746_ _0615_ _0884_ ZI_sky130_fd_sc_hd__a221o_2
X_8203_ VPWR VGND VGND VPWR _3572_ _3573_ _3571_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_88_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_11_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6395_ VGND VPWR VGND VPWR _1853_ _1438_ _1361_ _1349_ _1432_ _1289_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_112_153 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_88_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5346_ VGND VPWR _0816_ _0161_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_112_197 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8134_ VGND VPWR _3510_ _2637_ _2732_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8065_ VGND VPWR _3448_ _0365_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5277_ VGND VPWR _0747_ _0746_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7016_ VGND VPWR VGND VPWR _2468_ _2150_ _2194_ _2112_ ZI_sky130_fd_sc_hd__o21a_2
X_4228_ VPWR VGND VGND VPWR _3771_ _3762_ sword_ctr_reg\[1\] ZI_sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_106_Right_106 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7918_ VGND VPWR _3314_ _3311_ _3313_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7849_ VGND VPWR _3252_ _2549_ _3251_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_415 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_80_305 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_18_295 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_33_243 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_17_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_33_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_68_184 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_37_571 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_3_148 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_110_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6180_ VGND VPWR VGND VPWR _1641_ _1639_ _1453_ _1640_ _1432_ ZI_sky130_fd_sc_hd__a211o_2
X_5200_ VPWR VGND _0600_ _0670_ _0639_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_110_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5131_ VPWR VGND _0598_ _0601_ _0600_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5062_ VGND VPWR _0532_ _0531_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_74_76 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_74_54 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5964_ VGND VPWR _1426_ _1425_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7703_ VPWR VGND _3120_ block[93] round_key[93] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_90_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_75_600 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5895_ VGND VPWR VGND VPWR _1305_ _1333_ _1357_ _3850_ ZI_sky130_fd_sc_hd__a21oi_2
X_4915_ VGND VPWR _0389_ _0379_ _0388_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_97 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_7_410 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7634_ VGND VPWR _3056_ _4062_ _3055_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4846_ VGND VPWR VGND VPWR _4104_ new_block[99] _0320_ _0317_ _0294_ _0014_ ZI_sky130_fd_sc_hd__o32a_2
X_7565_ VGND VPWR VGND VPWR _2993_ _2992_ _2991_ _2989_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_74_176 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6516_ VPWR VGND VPWR VGND _1965_ _1971_ _1968_ _1787_ _1972_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_99_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4777_ VGND VPWR VGND VPWR _4104_ new_block[98] _0252_ _0247_ _0229_ _0013_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_43_585 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7496_ VGND VPWR _2930_ _2928_ _2929_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_602 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6447_ VGND VPWR VGND VPWR _1904_ _1893_ _1905_ _1001_ ZI_sky130_fd_sc_hd__a21oi_2
X_6378_ VGND VPWR _1837_ _1830_ _1836_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5329_ VGND VPWR _0799_ new_block[47] round_key[47] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8117_ VGND VPWR _3495_ _3493_ _3494_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8048_ VGND VPWR VGND VPWR _3331_ new_block[61] _3432_ _3429_ _2686_ _0104_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_65_198 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_110_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_104_473 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_88_246 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_56_132 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5680_ VPWR VGND _1146_ new_block[108] round_key[108] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_44_305 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4700_ VPWR VGND VGND VPWR _3992_ _0176_ _3859_ ZI_sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_7_Left_120 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_72_625 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4631_ _3803_ _4168_ _3794_ _3868_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7350_ VGND VPWR VGND VPWR _2796_ _4099_ _3770_ _3777_ ZI_sky130_fd_sc_hd__o21a_2
X_4562_ VGND VPWR VGND VPWR _4100_ _4099_ _4097_ _3777_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_12_246 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_40_533 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7281_ VPWR VGND VPWR VGND _2393_ _2728_ _2727_ _2358_ _2729_ ZI_sky130_fd_sc_hd__or4_2
X_6301_ VPWR VGND _1761_ _1760_ _1759_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4493_ VPWR VGND VGND VPWR _3929_ _4031_ _3803_ ZI_sky130_fd_sc_hd__nor2_2
X_6232_ VGND VPWR VGND VPWR _1693_ _1692_ _1691_ _1687_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_0_641 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6163_ VPWR VGND VGND VPWR _1549_ _1624_ _1495_ ZI_sky130_fd_sc_hd__nor2_2
X_6094_ VGND VPWR VGND VPWR _1555_ _1515_ _1474_ _1440_ _1556_ ZI_sky130_fd_sc_hd__a31o_2
X_5114_ VGND VPWR VGND VPWR _0583_ _0582_ _0584_ _0580_ _0577_ ZI_sky130_fd_sc_hd__nand4_2
X_5045_ VGND VPWR _0516_ _0514_ _0515_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_109_93 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_26_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6996_ VPWR VGND VPWR VGND _2285_ _2158_ _2208_ _2236_ _2448_ ZI_sky130_fd_sc_hd__a22o_2
X_5947_ _1319_ _1409_ _1353_ _1377_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_94_249 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5878_ VGND VPWR _1340_ _1339_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7617_ VPWR VGND _3041_ block[118] round_key[118] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4829_ VPWR VGND _0304_ _0303_ _0297_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_16_585 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7548_ VGND VPWR VGND VPWR _2894_ new_block[80] _2977_ _2975_ _1562_ _0059_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_16_596 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7479_ VPWR VGND _2914_ _1677_ _1568_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_39_611 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_30_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_93_293 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_111_218 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_39_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6850_ VGND VPWR VGND VPWR _2304_ _2299_ _2187_ _2301_ _2303_ ZI_sky130_fd_sc_hd__a211o_2
XPHY_EDGE_ROW_8_Right_8 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6781_ VPWR VGND _2105_ _2235_ _2129_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5801_ VGND VPWR VGND VPWR _1264_ _0610_ _0704_ _1262_ _1263_ ZI_sky130_fd_sc_hd__a211o_2
X_5732_ VPWR VGND _1197_ block[45] round_key[45] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8520_ VGND VPWR VPWR VGND clk _0122_ reset_n new_block[15] ZI_sky130_fd_sc_hd__dfrtp_2
X_5663_ VGND VPWR _1129_ _0998_ _1128_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8451_ VGND VPWR VPWR VGND clk _0053_ reset_n new_block[74] ZI_sky130_fd_sc_hd__dfrtp_2
X_5594_ VGND VPWR _1061_ _0799_ _0904_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_500 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8382_ VGND VPWR _3734_ _3731_ _3733_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4614_ VPWR VGND VPWR VGND _4151_ _4046_ ZI_sky130_fd_sc_hd__inv_2
X_7402_ VPWR VGND VPWR VGND _2797_ _2786_ _2843_ _2703_ _0431_ _2844_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_40_330 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4545_ VPWR VGND VGND VPWR _3760_ _4083_ dec_ctrl_reg\[1\] ZI_sky130_fd_sc_hd__nor2_2
X_7333_ VPWR VGND _2780_ _0523_ _0363_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4476_ VPWR VGND VPWR VGND _4013_ _3950_ _3911_ _4012_ _4014_ ZI_sky130_fd_sc_hd__a22o_2
X_7264_ VGND VPWR VGND VPWR _2712_ _2222_ _2155_ _2144_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_96_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6215_ VPWR VGND _1676_ round_key[16] new_block[16] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_39_Right_39 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7195_ VPWR VGND _2645_ block[124] round_key[124] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_96_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6146_ VPWR VGND VPWR VGND _1603_ _1606_ _1605_ _1602_ _1607_ ZI_sky130_fd_sc_hd__or4_2
X_6077_ VPWR VGND VGND VPWR _1416_ _1539_ _1538_ ZI_sky130_fd_sc_hd__nor2_2
X_5028_ VPWR VGND VGND VPWR _3955_ _0499_ _3954_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_67_205 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6979_ VPWR VGND VPWR VGND _2373_ _2216_ _2102_ _2144_ _2431_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_35_113 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_36_625 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_106_502 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_50_105 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_63_477 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Right_57 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_25_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Left_201 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Right_66 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_58_227 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_81_241 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_42_628 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_54_477 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_112_505 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_81_296 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_54_499 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_34_190 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_97_Left_210 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Right_75 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4330_ VPWR VGND VGND VPWR _3775_ _3868_ _3814_ _3809_ ZI_sky130_fd_sc_hd__nor3b_2
X_4261_ VGND VPWR VGND VPWR _3799_ new_block[33] sword_ctr_reg\[1\] sword_ctr_reg\[0\]
+ ZI_sky130_fd_sc_hd__and3b_2
XFILLER_0_5_69 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6000_ VGND VPWR _1462_ _1461_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7951_ VPWR VGND _3344_ _0380_ _0373_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_84_Right_84 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7882_ VGND VPWR _3282_ _3280_ _3281_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6902_ VPWR VGND _2118_ _2355_ _2162_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_82_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6833_ VPWR VGND VPWR VGND _2286_ _2230_ _2223_ _2136_ _2171_ _2287_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_9_302 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_106_94 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_92_517 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_9_346 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_17_102 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6764_ _2070_ _2218_ _2182_ _2162_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8503_ VGND VPWR VPWR VGND clk _0105_ reset_n new_block[62] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_455 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5715_ VPWR VGND VPWR VGND _1174_ _1179_ _1176_ _1167_ _1180_ ZI_sky130_fd_sc_hd__or4_2
X_6695_ VGND VPWR _2149_ _2148_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_31_80 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_33_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5646_ VGND VPWR VGND VPWR _1112_ _0734_ _0545_ _0888_ _0709_ _0589_ ZI_sky130_fd_sc_hd__a32o_2
X_8434_ VGND VPWR VPWR VGND clk _0036_ reset_n new_block[121] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_60_414 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_93_Right_93 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_72_296 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5577_ VPWR VGND VPWR VGND _1044_ _1042_ _1043_ ZI_sky130_fd_sc_hd__or2_2
X_8365_ VPWR VGND VGND VPWR _3719_ _1897_ _3718_ ZI_sky130_fd_sc_hd__nand2_2
X_8296_ VPWR VGND _3657_ block[53] round_key[53] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7316_ VPWR VGND VPWR VGND _2601_ _2762_ _2759_ _2251_ _2763_ ZI_sky130_fd_sc_hd__or4_2
X_4528_ VGND VPWR _4066_ new_block[71] round_key[71] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_193 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7247_ VGND VPWR _2696_ _2315_ _2695_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4459_ VPWR VGND VGND VPWR _3877_ _3997_ _3803_ ZI_sky130_fd_sc_hd__nor2_2
X_7178_ VGND VPWR _2628_ _1961_ _2409_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6129_ VPWR VGND VGND VPWR _1524_ _1590_ _1447_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_99_105 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_95_388 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_55_219 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_36_433 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_36_444 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_24_639 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_36_499 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_51_425 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_15_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5500_ VGND VPWR VPWR VGND _0966_ _0967_ _0611_ _0968_ ZI_sky130_fd_sc_hd__or3_2
X_6480_ VPWR VGND VPWR VGND _1931_ _1936_ _1933_ _1784_ _1937_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_2_533 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5431_ VPWR VGND _0900_ round_key[57] new_block[57] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8150_ VPWR VGND _3525_ _2048_ _0489_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5362_ VPWR VGND VPWR VGND _0718_ _0602_ _0740_ _0619_ _0706_ _0831_ ZI_sky130_fd_sc_hd__a221o_2
X_7101_ VGND VPWR _2552_ _0920_ _1241_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4313_ VGND VPWR VGND VPWR _3814_ _3809_ _3851_ _3850_ ZI_sky130_fd_sc_hd__a21oi_2
X_8081_ VGND VPWR VGND VPWR _3462_ new_block[0] _3460_ _3456_ _4060_ _0107_ ZI_sky130_fd_sc_hd__o32a_2
X_5293_ VPWR VGND _0600_ _0763_ _0596_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_7032_ VGND VPWR _2484_ _0250_ _0523_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4244_ VGND VPWR VGND VPWR _3782_ round[2] _3784_ _0000_ ZI_sky130_fd_sc_hd__a21oi_2
X_7934_ VPWR VGND _3329_ block[83] round_key[83] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7865_ VPWR VGND _3267_ block[108] round_key[108] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6816_ VGND VPWR VPWR VGND _2268_ _2269_ _2266_ _2270_ ZI_sky130_fd_sc_hd__or3_2
X_7796_ VGND VPWR _3204_ _1828_ _1945_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_517 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6747_ VGND VPWR _2201_ _2200_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6678_ VGND VPWR _2132_ _2131_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_73_583 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8417_ VGND VPWR VPWR VGND clk _0019_ reset_n new_block[104] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_233 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5629_ VGND VPWR VGND VPWR _1095_ _0729_ _0635_ _0661_ _0671_ _0674_ ZI_sky130_fd_sc_hd__a32o_2
X_8348_ VPWR VGND _3704_ block[26] round_key[26] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8279_ VGND VPWR _3641_ _1069_ _1139_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_68_344 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_56_506 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_28_208 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_107_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_32_491 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_129 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5980_ _1295_ _1442_ _1400_ _1441_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_59_322 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4931_ VPWR VGND VGND VPWR _3862_ _3849_ _0404_ _4016_ _3975_ ZI_sky130_fd_sc_hd__o22ai_2
XFILLER_0_87_642 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4862_ VGND VPWR VGND VPWR _3969_ _4036_ _3988_ _3999_ _0336_ ZI_sky130_fd_sc_hd__o22a_2
X_7650_ VPWR VGND _3071_ block[89] round_key[89] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_86_174 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_74_347 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6601_ VGND VPWR VGND VPWR _2055_ new_block[60] sword_ctr_reg\[1\] sword_ctr_reg\[0\]
+ ZI_sky130_fd_sc_hd__and3b_2
X_7581_ VGND VPWR VGND VPWR _2997_ new_block[83] _3007_ _3005_ _1815_ _0062_ ZI_sky130_fd_sc_hd__o32a_2
XPHY_EDGE_ROW_25_Left_138 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_103_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_62_509 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_55_561 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4793_ VGND VPWR VGND VPWR _3987_ _4115_ _3955_ _4052_ _0268_ ZI_sky130_fd_sc_hd__o22a_2
X_6532_ _1308_ _1988_ _1424_ _1409_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_42_200 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6463_ VGND VPWR VGND VPWR _1542_ _1336_ _1917_ _1918_ _1920_ _1919_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_30_406 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5414_ VGND VPWR VGND VPWR _0883_ _0626_ _0705_ _0583_ _0630_ ZI_sky130_fd_sc_hd__and4_2
X_8202_ VGND VPWR VGND VPWR _3570_ _3569_ _0158_ _3572_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_88_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6394_ VPWR VGND VPWR VGND _1852_ _1789_ _1851_ ZI_sky130_fd_sc_hd__or2_2
XFILLER_0_112_165 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_88_97 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8133_ VGND VPWR VGND VPWR _3462_ new_block[5] _3509_ _3507_ _0429_ _0112_ ZI_sky130_fd_sc_hd__o32a_2
X_5345_ VGND VPWR VPWR VGND _0813_ _0804_ _0815_ _0444_ _0814_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_10_141 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8064_ VPWR VGND VGND VPWR _3447_ _3445_ _3446_ ZI_sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_34_Left_147 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5276_ VGND VPWR _0746_ _0745_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7015_ VGND VPWR VGND VPWR _2219_ _2465_ _2381_ _2466_ _2467_ ZI_sky130_fd_sc_hd__o22a_2
X_4227_ VPWR VGND VGND VPWR _3770_ sword_ctr_reg\[0\] _3764_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_37_90 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7917_ VGND VPWR _3313_ _3134_ _3312_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_38_517 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Left_156 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_93_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7848_ VGND VPWR _3251_ _2978_ _3250_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7779_ VGND VPWR VGND VPWR _3153_ new_block[36] _3188_ _3186_ _0362_ _0079_ ZI_sky130_fd_sc_hd__o32a_2
XPHY_EDGE_ROW_52_Left_165 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_17_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_108_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_174 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_29_517 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_84_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_37_583 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_83_188 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_71_328 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_3_105 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_70_Left_183 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_110_625 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5130_ VGND VPWR _0600_ _0599_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5061_ VPWR VGND VGND VPWR _0531_ _3754_ _0530_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_74_66 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5963_ _1362_ _1425_ _1352_ _1413_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_4914_ VGND VPWR _0388_ _0381_ _0387_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7702_ VGND VPWR VPWR VGND _3116_ _3115_ _3119_ _3118_ _3117_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_75_612 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5894_ VGND VPWR VGND VPWR _1356_ _1355_ _1351_ _1346_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_90_65 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_47_369 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7633_ VGND VPWR _3055_ _4061_ _0142_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_615 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4845_ VPWR VGND VPWR VGND _4101_ _0169_ _0319_ _0162_ _0318_ _0320_ ZI_sky130_fd_sc_hd__a221o_2
X_7564_ VGND VPWR VGND VPWR _2991_ _2989_ _2992_ _2642_ ZI_sky130_fd_sc_hd__a21oi_2
X_4776_ VGND VPWR VGND VPWR _0251_ _4094_ _0248_ _0249_ _0252_ ZI_sky130_fd_sc_hd__a31o_2
X_6515_ VGND VPWR VGND VPWR _1434_ _1308_ _1492_ _1969_ _1971_ _1970_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_15_288 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_43_597 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7495_ VGND VPWR _2929_ _1888_ _1901_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6446_ VGND VPWR _1904_ _1894_ _1903_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_124 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6377_ VGND VPWR _1836_ _1831_ _1835_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5328_ VPWR VGND _0798_ _0797_ _0794_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8116_ VGND VPWR _3494_ _2631_ _3011_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8047_ VGND VPWR VGND VPWR _3432_ _3430_ _2857_ _3431_ _3150_ ZI_sky130_fd_sc_hd__a211o_2
X_5259_ VGND VPWR _0729_ _0728_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_97_269 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_78_472 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_66_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_93_420 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_66_645 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_19_550 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_28_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_57_601 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4630_ VGND VPWR VGND VPWR _4166_ _4165_ _4167_ _4164_ _4163_ ZI_sky130_fd_sc_hd__nand4_2
XFILLER_0_52_361 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4561_ VGND VPWR _4099_ _4098_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_71_169 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6300_ VPWR VGND _1760_ _1676_ _1570_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_8_69 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7280_ VPWR VGND VPWR VGND _2338_ _2155_ _2336_ _2214_ _2728_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_69_44 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4492_ _3838_ _4030_ _3890_ _3901_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_100_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6231_ VGND VPWR VGND VPWR _1691_ _1687_ _1692_ _1001_ ZI_sky130_fd_sc_hd__a21oi_2
X_6162_ VPWR VGND VPWR VGND _1596_ _1622_ _1612_ _1374_ _1623_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_40_589 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5113_ VGND VPWR _0583_ _0557_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_110_477 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6093_ _1424_ _1555_ _1394_ _1361_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5044_ VPWR VGND _0515_ _0373_ _0142_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_108_Left_221 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_19_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_79_247 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6995_ _2205_ _2447_ _2126_ _2157_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5946_ VGND VPWR _1408_ _1407_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_48_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5877_ _1312_ _1339_ _1338_ _1318_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7616_ VGND VPWR VPWR VGND _3038_ _3037_ _3040_ _2855_ _3039_ ZI_sky130_fd_sc_hd__o211a_2
X_4828_ VGND VPWR _0303_ _0299_ _0302_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_626 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_47_199 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_90_456 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_62_158 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_62_136 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7547_ VPWR VGND VPWR VGND _2892_ _2976_ _2857_ _2880_ _4075_ _2977_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_31_501 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4759_ VGND VPWR _0235_ _4075_ _4073_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_372 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7478_ VGND VPWR _2913_ _1835_ _2912_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6429_ VGND VPWR _1887_ _1885_ _1886_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_109_500 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_93_261 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_34_361 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_22_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_55_57 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_55_46 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_29_100 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6780_ VPWR VGND _2170_ _2234_ _2184_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_71_45 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5800_ VGND VPWR VGND VPWR _1263_ _0628_ _0546_ _0619_ _0775_ _0923_ ZI_sky130_fd_sc_hd__a32o_2
X_5731_ VGND VPWR VGND VPWR _1196_ _1195_ _1194_ _1191_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_57_486 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5662_ VPWR VGND _1128_ _1072_ _0802_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8450_ VGND VPWR VPWR VGND clk _0052_ reset_n new_block[73] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_72_456 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5593_ VGND VPWR _1060_ _0986_ _1059_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_309 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8381_ VGND VPWR _3733_ _2039_ _3732_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7401_ VPWR VGND _2843_ block[36] round_key[36] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4613_ VGND VPWR VGND VPWR _4150_ _3913_ _3881_ _4148_ _4149_ ZI_sky130_fd_sc_hd__a211o_2
X_7332_ VGND VPWR _2779_ _2776_ _2778_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_52_180 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_111_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4544_ VPWR VGND VPWR VGND _4082_ _3772_ _3767_ ZI_sky130_fd_sc_hd__or2_2
X_7263_ VGND VPWR VGND VPWR _2711_ _2709_ _2132_ _2710_ _2465_ ZI_sky130_fd_sc_hd__a211o_2
X_6214_ VGND VPWR VPWR VGND _1675_ _1623_ _1643_ _1674_ _3755_ ZI_sky130_fd_sc_hd__o31a_2
X_4475_ _3878_ _4013_ _3794_ _3815_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_96_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7194_ VGND VPWR VGND VPWR _2644_ _2643_ _2641_ _2636_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_110_263 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6145_ VPWR VGND VGND VPWR _1466_ _1606_ _1401_ ZI_sky130_fd_sc_hd__nor2_2
X_6076_ VGND VPWR _1538_ _1537_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5027_ VGND VPWR VGND VPWR _3926_ _4189_ _4047_ _4135_ _0498_ _4171_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_67_217 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6978_ VGND VPWR VGND VPWR _2185_ _2343_ _2372_ _2230_ _2430_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_0_81 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5929_ VPWR VGND VGND VPWR _1391_ _3754_ _1300_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_36_637 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_48_486 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_75_250 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_106_514 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_63_456 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_63_489 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_39_464 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_39_475 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_26_125 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_14_309 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_54_489 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_81_286 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_112_517 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4260_ sword_ctr_reg\[1\] _3798_ sword_ctr_reg\[0\] new_block[1] VPWR VGND VPWR VGND
+ ZI_sky130_fd_sc_hd__and3_2
X_7950_ VGND VPWR VGND VPWR _3331_ new_block[52] _3343_ _3341_ _1884_ _0095_ ZI_sky130_fd_sc_hd__o32a_2
X_6901_ VGND VPWR VGND VPWR _2354_ _2255_ _2227_ _2173_ ZI_sky130_fd_sc_hd__o21a_2
X_7881_ VPWR VGND _3281_ _2733_ _0447_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6832_ VPWR VGND VPWR VGND _2255_ _2285_ _2135_ _2144_ _2286_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_82_99 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6763_ VPWR VGND _2184_ _2217_ _2216_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_57_250 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8502_ VGND VPWR VPWR VGND clk _0104_ reset_n new_block[61] ZI_sky130_fd_sc_hd__dfrtp_2
X_5714_ VPWR VGND VPWR VGND _0736_ _0768_ _1179_ _0699_ _1178_ ZI_sky130_fd_sc_hd__or4b_2
X_6694_ VPWR VGND VGND VPWR _2147_ _2148_ _2146_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_72_220 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_33_629 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8433_ VGND VPWR VPWR VGND clk _0035_ reset_n new_block[120] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_489 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5645_ _0612_ _1111_ _0688_ _0841_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_72_253 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_86_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5576_ VPWR VGND VPWR VGND _0785_ _0692_ _0645_ _0666_ _1043_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_41_662 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8364_ VGND VPWR _3718_ _2930_ _3717_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_386 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8295_ VGND VPWR VPWR VGND _3654_ _2833_ _3656_ _0366_ _3655_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_40_161 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4527_ VPWR VGND _4065_ _4064_ _4061_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7315_ VPWR VGND VPWR VGND _2372_ _2761_ _2327_ _2171_ _2762_ ZI_sky130_fd_sc_hd__a22o_2
X_7246_ VGND VPWR _2695_ _1055_ _1280_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_561 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4458_ VPWR VGND VPWR VGND _3986_ _3995_ _3996_ _3981_ _3985_ ZI_sky130_fd_sc_hd__or4b_2
X_7177_ VGND VPWR _2627_ _2625_ _2626_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6128_ VPWR VGND VPWR VGND _1588_ _1531_ _1444_ _1426_ _1589_ ZI_sky130_fd_sc_hd__a22o_2
X_4389_ VPWR VGND VPWR VGND _3926_ _3925_ _3913_ _3923_ _3927_ ZI_sky130_fd_sc_hd__a22o_2
X_6059_ VGND VPWR _1521_ _1289_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_68_515 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_36_456 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_106_300 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_106_322 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_31_150 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_36_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_67_570 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_54_220 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_6_339 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_54_253 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_15_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5430_ VGND VPWR VGND VPWR _0899_ _3756_ _0898_ _0832_ ZI_sky130_fd_sc_hd__o21a_2
X_5361_ VGND VPWR VGND VPWR _0830_ _0825_ _0669_ _0826_ _0829_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_2_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_10_323 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7100_ VGND VPWR _2551_ _1055_ _2550_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5292_ VGND VPWR VGND VPWR _0762_ _0678_ _0696_ _0602_ ZI_sky130_fd_sc_hd__o21a_2
X_8080_ VGND VPWR _3462_ _3461_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4312_ VGND VPWR _3850_ _3832_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7031_ VGND VPWR VPWR VGND _2471_ _2482_ _2460_ _2483_ ZI_sky130_fd_sc_hd__or3_2
X_4243_ VGND VPWR _0008_ _3783_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7933_ VGND VPWR _3328_ _2702_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_89_183 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7864_ VGND VPWR VPWR VGND _3263_ _3259_ _3266_ _3265_ _3264_ ZI_sky130_fd_sc_hd__o211a_2
X_6815_ VPWR VGND _2096_ _2269_ _2184_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_7795_ VGND VPWR _3203_ _1950_ _3202_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_529 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_42_80 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6746_ VPWR VGND _2199_ _2200_ _2105_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_9_177 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6677_ VGND VPWR _2131_ _2130_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5628_ VPWR VGND VPWR VGND _0620_ _0834_ _0746_ _0678_ _1094_ ZI_sky130_fd_sc_hd__a22o_2
X_8416_ VGND VPWR VPWR VGND clk _0018_ reset_n new_block[103] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_109 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8347_ VGND VPWR VPWR VGND _3701_ _3700_ _3703_ _0366_ _3702_ ZI_sky130_fd_sc_hd__o211a_2
X_5559_ VGND VPWR VGND VPWR _1026_ _0651_ _0740_ _0589_ ZI_sky130_fd_sc_hd__o21a_2
X_8278_ VGND VPWR VGND VPWR _3640_ new_block[19] _3639_ _3637_ _1815_ _0126_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_6_80 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7229_ VPWR VGND VPWR VGND _2672_ _2677_ _2674_ _2254_ _2678_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_95_142 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_83_304 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_107_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_91_381 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_102_391 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_87_610 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_63_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_87_654 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4930_ VGND VPWR VGND VPWR _0399_ _3920_ _0401_ _0402_ _0403_ _0323_ ZI_sky130_fd_sc_hd__a2111o_2
X_4861_ VGND VPWR VGND VPWR _3987_ _4021_ _3872_ _3988_ _0335_ ZI_sky130_fd_sc_hd__o22a_2
XFILLER_0_86_164 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_86_186 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6600_ VGND VPWR VGND VPWR _3797_ _2050_ _2051_ _2052_ _2054_ _2053_ ZI_sky130_fd_sc_hd__o41ai_2
X_7580_ VPWR VGND VPWR VGND _2995_ _2960_ _3006_ _2984_ _0308_ _3007_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_74_359 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4792_ VGND VPWR VGND VPWR _0267_ _4031_ _3925_ _0265_ _0266_ ZI_sky130_fd_sc_hd__a211o_2
X_6531_ VPWR VGND _1499_ _1987_ _1443_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_27_264 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_42_212 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_103_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_6_169 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6462_ VGND VPWR VGND VPWR _1464_ _1557_ _1660_ _1670_ _1919_ _1742_ ZI_sky130_fd_sc_hd__a2111o_2
X_6393_ VPWR VGND VPWR VGND _1811_ _1603_ _1525_ _1422_ _1851_ ZI_sky130_fd_sc_hd__or4_2
X_5413_ VGND VPWR VPWR VGND _0879_ _0881_ _0878_ _0882_ ZI_sky130_fd_sc_hd__or3_2
X_8201_ VPWR VGND VGND VPWR _3570_ _3571_ _3569_ ZI_sky130_fd_sc_hd__nor2_2
X_5344_ VPWR VGND VGND VPWR _0814_ _0804_ _0813_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_88_65 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8132_ VPWR VGND VPWR VGND _3459_ _3490_ _3508_ _3468_ _1564_ _3509_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_10_153 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_11_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8063_ VPWR VGND _3446_ _2867_ _2849_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5275_ VPWR VGND _0598_ _0745_ _0578_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_10_197 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7014_ VGND VPWR VGND VPWR _2159_ _2228_ _2127_ _2466_ ZI_sky130_fd_sc_hd__a21o_2
X_4226_ VGND VPWR _0005_ _3769_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7916_ VGND VPWR _3312_ _4075_ _0154_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7847_ VPWR VGND _3250_ _2639_ _2565_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_93_613 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_65_337 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_46_551 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_92_167 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7778_ VPWR VGND VPWR VGND _3150_ _3159_ _3187_ _3139_ _1132_ _3188_ ZI_sky130_fd_sc_hd__a221o_2
X_6729_ VPWR VGND _2182_ _2183_ _2139_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_104_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_104_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_84_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_68_197 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_56_348 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_110_637 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_20_473 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5060_ VGND VPWR VPWR VGND _0528_ _0527_ _0526_ _3828_ _0529_ _0530_ ZI_sky130_fd_sc_hd__a41oi_2
X_5962_ VGND VPWR _1424_ _1400_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4913_ VGND VPWR _0387_ _0384_ _0386_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_87_462 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7701_ VGND VPWR _3118_ _0365_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5893_ VGND VPWR _1355_ _1354_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_90_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_74_112 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7632_ VGND VPWR _3054_ _4075_ _0150_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_134 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4844_ VPWR VGND _0319_ round_key[99] new_block[99] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7563_ VGND VPWR _2991_ _2633_ _2990_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_627 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4775_ VGND VPWR _4103_ _4090_ _0251_ _0250_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
X_6514_ VPWR VGND VPWR VGND _1359_ _1616_ _1308_ _1511_ _1970_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_43_543 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7494_ VGND VPWR _2928_ _1682_ _1765_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_215 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6445_ VGND VPWR _1903_ _1897_ _1902_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6376_ VGND VPWR _1835_ _1832_ _1834_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5327_ VPWR VGND _0797_ _0796_ _0795_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8115_ VGND VPWR _3493_ _1908_ _3492_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8046_ VPWR VGND VGND VPWR _0805_ _3431_ _4090_ ZI_sky130_fd_sc_hd__nor2_2
X_5258_ VPWR VGND VGND VPWR _0649_ _0728_ _0629_ ZI_sky130_fd_sc_hd__nor2_2
X_5189_ VGND VPWR VGND VPWR _0659_ _0656_ _0655_ _0571_ _0658_ _0654_ ZI_sky130_fd_sc_hd__a32o_2
X_4209_ sword_ctr_reg\[1\] _3757_ sword_ctr_reg\[0\] dec_ctrl_reg\[1\] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_3_81 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_97_204 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_66_613 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_65_189 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_80_148 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_21_204 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_0_109 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_61_384 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_69_440 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_84_421 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4560_ VPWR VGND _4089_ _4098_ _4082_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_8_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_25_554 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_25_576 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_107_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4491_ _3924_ _4029_ _3881_ _3939_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_100_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6230_ VGND VPWR _1691_ _1581_ _1690_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6161_ VPWR VGND VPWR VGND _1618_ _1621_ _1620_ _1615_ _1622_ ZI_sky130_fd_sc_hd__or4_2
X_5112_ VGND VPWR _0582_ _0581_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_110_489 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6092_ VGND VPWR VGND VPWR _1376_ _1340_ _1546_ _1550_ _1554_ _1553_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_85_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5043_ VGND VPWR _0514_ _0230_ _0376_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_109_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_48_602 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6994_ VPWR VGND VPWR VGND _2441_ _2445_ _2442_ _2439_ _2446_ ZI_sky130_fd_sc_hd__or4_2
X_5945_ _1335_ _1407_ _1334_ _1295_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_87_281 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5876_ VPWR VGND VGND VPWR _3775_ _1324_ _1329_ _1338_ ZI_sky130_fd_sc_hd__nor3_2
XFILLER_0_48_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7615_ VPWR VGND VGND VPWR _3039_ _3037_ _3038_ ZI_sky130_fd_sc_hd__nand2_2
X_4827_ VPWR VGND _0302_ _0301_ _4064_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_63_649 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4758_ VPWR VGND _0234_ round_key[82] new_block[82] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7546_ VPWR VGND _2976_ block[112] round_key[112] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_31_513 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7477_ VPWR VGND _2912_ _1891_ _1819_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4689_ VPWR VGND VPWR VGND _0166_ dec_ctrl_reg\[2\] ZI_sky130_fd_sc_hd__inv_2
XFILLER_0_31_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6428_ VGND VPWR _1886_ _1570_ _1821_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_445 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_11_281 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6359_ VGND VPWR _1818_ _1580_ _1817_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8029_ VPWR VGND _3415_ _3414_ _1188_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_14_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_39_624 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_38_156 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_93_273 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_53_159 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5730_ VGND VPWR VGND VPWR _1194_ _1191_ _1195_ _1001_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_71_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_84_273 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5661_ VPWR VGND _1127_ _1126_ _0914_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7400_ VPWR VGND VGND VPWR _2841_ _2842_ _0158_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_57_498 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5592_ VPWR VGND _1059_ _1058_ _0797_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4612_ VPWR VGND VGND VPWR _4116_ _4110_ _4149_ _4114_ _4121_ ZI_sky130_fd_sc_hd__o22ai_2
X_8380_ VPWR VGND _3732_ _1819_ _1574_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7331_ VGND VPWR _2778_ _2411_ _2777_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4543_ VPWR VGND VGND VPWR _4080_ _4081_ _4071_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_13_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_52_192 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7262_ VGND VPWR VGND VPWR _2710_ _2259_ _2203_ _2187_ _2373_ _2207_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_102_209 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6213_ VPWR VGND VPWR VGND _1666_ _1673_ _1669_ _1659_ _1674_ ZI_sky130_fd_sc_hd__or4_2
X_4474_ _3838_ _4012_ _3831_ _3892_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7193_ VGND VPWR VGND VPWR _2641_ _2636_ _2643_ _2642_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_110_253 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_96_65 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6144_ _1414_ _1605_ _1319_ _1604_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_96_98 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6075_ VGND VPWR VPWR VGND _1393_ _1455_ _1391_ _1537_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_31_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5026_ VPWR VGND VPWR VGND _4032_ _0205_ _0200_ _4006_ _0497_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_48_421 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6977_ VPWR VGND VPWR VGND _2426_ _2428_ _2427_ _2425_ _2429_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_95_549 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5928_ VGND VPWR _1390_ _1389_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_63_413 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5859_ VGND VPWR VGND VPWR _1321_ new_block[53] sword_ctr_reg\[1\] sword_ctr_reg\[0\]
+ ZI_sky130_fd_sc_hd__and3b_2
XFILLER_0_48_498 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_106_526 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7529_ VPWR VGND VPWR VGND _2892_ _2960_ _2959_ _2880_ _0153_ _2961_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_43_181 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_101_220 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_25_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_41_16 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_81_276 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_112_529 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_10_516 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_5_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_66_68 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7880_ VGND VPWR _3280_ _2689_ _3279_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6900_ VPWR VGND VPWR VGND _2186_ _2157_ _2096_ _2195_ _2353_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_106_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6831_ VGND VPWR _2285_ _2201_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6762_ VGND VPWR _2216_ _2215_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8501_ VGND VPWR VPWR VGND clk _0103_ reset_n new_block[60] ZI_sky130_fd_sc_hd__dfrtp_2
X_5713_ VPWR VGND VPWR VGND _1177_ _0747_ _0740_ _0706_ _0689_ _1178_ ZI_sky130_fd_sc_hd__a221o_2
X_6693_ VGND VPWR VPWR VGND _2104_ _2083_ _3775_ _2147_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_72_232 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_26_660 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8432_ VGND VPWR VPWR VGND clk _0034_ reset_n new_block[119] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_468 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5644_ VGND VPWR VGND VPWR _1110_ _0710_ _0757_ _1107_ _1109_ ZI_sky130_fd_sc_hd__a211o_2
X_8363_ VGND VPWR _3717_ _2007_ _3716_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_587 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5575_ VGND VPWR VGND VPWR _1042_ _0746_ _0712_ _0645_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_103_518 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7314_ VPWR VGND VPWR VGND _2761_ _2178_ _2760_ ZI_sky130_fd_sc_hd__or2_2
X_8294_ VPWR VGND VGND VPWR _3655_ _2833_ _3654_ ZI_sky130_fd_sc_hd__nand2_2
X_4526_ VGND VPWR _4064_ _4062_ _4063_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_173 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7245_ VPWR VGND _2694_ _2646_ _1908_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4457_ VPWR VGND VGND VPWR _3988_ _3933_ _3987_ _3974_ _3995_ _3994_ ZI_sky130_fd_sc_hd__o221a_2
XFILLER_0_0_281 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7176_ VGND VPWR _2626_ _1908_ _2547_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6127_ VPWR VGND VGND VPWR _1307_ _1588_ _1336_ ZI_sky130_fd_sc_hd__nor2_2
X_4388_ VPWR VGND _3815_ _3926_ _3920_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_6058_ VPWR VGND VPWR VGND _1519_ _1518_ _1397_ _1345_ _1379_ _1520_ ZI_sky130_fd_sc_hd__a221o_2
X_5009_ VGND VPWR _0481_ _0480_ _0432_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_313 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_68_527 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_63_232 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_51_449 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_31_162 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_99_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Right_101 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_59_505 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_52_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_86_357 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_109_150 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_54_232 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_54_287 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_23_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5360_ VGND VPWR VGND VPWR _0828_ _0620_ _0827_ _0757_ _0829_ ZI_sky130_fd_sc_hd__a31o_2
X_5291_ _0592_ _0761_ _0557_ _0569_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_4311_ VGND VPWR _3849_ _3848_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7030_ VPWR VGND VPWR VGND _2476_ _2481_ _2477_ _2474_ _2482_ ZI_sky130_fd_sc_hd__or4_2
X_4242_ VPWR VGND VPWR VGND _3782_ _3783_ _0000_ _3781_ ZI_sky130_fd_sc_hd__or3b_2
X_7932_ VGND VPWR VPWR VGND _3325_ _3324_ _3327_ _3265_ _3326_ ZI_sky130_fd_sc_hd__o211a_2
X_7863_ VGND VPWR _3265_ _0365_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_89_195 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_92_316 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7794_ VGND VPWR _3202_ _1689_ _1817_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6814_ VGND VPWR VGND VPWR _2268_ _2267_ _2170_ _2106_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_45_221 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6745_ VGND VPWR VGND VPWR _2094_ _2089_ _3774_ _2199_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_58_582 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6676_ VPWR VGND _2128_ _2130_ _2129_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_8415_ VGND VPWR VPWR VGND clk _0017_ reset_n new_block[102] ZI_sky130_fd_sc_hd__dfrtp_2
X_5627_ VGND VPWR VGND VPWR _0740_ _0546_ _0854_ _1093_ ZI_sky130_fd_sc_hd__a21o_2
X_8346_ VPWR VGND VGND VPWR _3702_ _3700_ _3701_ ZI_sky130_fd_sc_hd__nand2_2
X_5558_ VPWR VGND VPWR VGND _1025_ _0736_ _0834_ ZI_sky130_fd_sc_hd__or2_2
XFILLER_0_41_482 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8277_ VGND VPWR _3640_ _3461_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4509_ VGND VPWR VGND VPWR _4047_ _3892_ _3868_ _3891_ _3890_ ZI_sky130_fd_sc_hd__and4_2
X_5489_ VPWR VGND VPWR VGND _0951_ _0956_ _0957_ _0694_ _0945_ ZI_sky130_fd_sc_hd__or4b_2
XFILLER_0_111_381 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7228_ VPWR VGND VGND VPWR _2676_ _2675_ _2099_ _2182_ _2336_ _2677_ ZI_sky130_fd_sc_hd__a311o_2
X_7159_ VGND VPWR VGND VPWR _2609_ _2138_ _2133_ _2105_ _2252_ ZI_sky130_fd_sc_hd__and4_2
XFILLER_0_95_154 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_107_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_106_197 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_20_611 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_86_110 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_63_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4860_ VPWR VGND VPWR VGND _0333_ _0334_ _0321_ _0324_ ZI_sky130_fd_sc_hd__or3b_2
XFILLER_0_87_666 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6530_ VPWR VGND VPWR VGND _1862_ _1986_ _1984_ _1985_ ZI_sky130_fd_sc_hd__or3b_2
X_4791_ VPWR VGND VGND VPWR _3976_ _0266_ _3851_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_55_541 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_12_73 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6461_ VGND VPWR VGND VPWR _1475_ _1655_ _1918_ _1549_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_42_224 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_103_97 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_70_533 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_11_600 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6392_ VPWR VGND VPWR VGND _1773_ _1849_ _1647_ _1615_ _1850_ ZI_sky130_fd_sc_hd__or4_2
X_5412_ VPWR VGND VPWR VGND _0880_ _0677_ _0825_ _0739_ _0751_ _0881_ ZI_sky130_fd_sc_hd__a221o_2
X_8200_ VPWR VGND _3570_ _3096_ _0368_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5343_ VGND VPWR _0813_ _0807_ _0812_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_110 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_88_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8131_ VPWR VGND _3508_ block[101] round_key[101] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8062_ VGND VPWR _3445_ _1272_ _3444_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_165 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5274_ VGND VPWR VGND VPWR _0744_ _0668_ _0657_ _0601_ ZI_sky130_fd_sc_hd__o21a_2
X_7013_ VPWR VGND _2345_ _2465_ _2355_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_4225_ VGND VPWR VPWR VGND sword_ctr_reg\[0\] _3768_ _3756_ _3769_ ZI_sky130_fd_sc_hd__mux2_2
XFILLER_0_97_419 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7915_ VGND VPWR _3311_ _0147_ _0430_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7846_ VGND VPWR VGND VPWR _3240_ new_block[42] _3249_ _3247_ _0984_ _0085_ ZI_sky130_fd_sc_hd__o32a_2
X_4989_ VPWR VGND VPWR VGND _0212_ _0266_ _0261_ _0191_ _0461_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_65_349 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7777_ VPWR VGND _3187_ block[4] round_key[4] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_46_585 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6728_ VGND VPWR _2182_ _2121_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_104_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6659_ VGND VPWR VGND VPWR _2113_ _2064_ _2063_ _2069_ _3753_ ZI_sky130_fd_sc_hd__and4_2
XFILLER_0_104_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8329_ VGND VPWR VGND VPWR _3640_ new_block[24] _3686_ _3684_ _2307_ _0131_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_68_110 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_33_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_68_165 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_68_132 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_56_305 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_83_113 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_37_530 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_52_533 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_52_599 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5961_ VGND VPWR VGND VPWR _1423_ _1355_ _1395_ _1417_ _1422_ ZI_sky130_fd_sc_hd__a211o_2
X_4912_ VGND VPWR _0386_ _0143_ _0385_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7700_ VPWR VGND VGND VPWR _3117_ _3115_ _3116_ ZI_sky130_fd_sc_hd__nand2_2
X_5892_ _1319_ _1354_ _1353_ _1330_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7631_ VGND VPWR VGND VPWR _2997_ new_block[87] _3053_ _3050_ _2038_ _0066_ ZI_sky130_fd_sc_hd__o32a_2
X_4843_ VPWR VGND _0318_ block[67] round_key[67] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_74_157 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7562_ VGND VPWR _2990_ _1586_ _2552_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_639 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4774_ VGND VPWR _0250_ new_block[98] round_key[98] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6513_ VPWR VGND VGND VPWR _1609_ _1969_ _1655_ ZI_sky130_fd_sc_hd__nor2_2
X_7493_ VGND VPWR _2927_ _2925_ _2926_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_382 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_43_555 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6444_ VGND VPWR _1902_ _1900_ _1901_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_30_227 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6375_ VGND VPWR _1834_ _1683_ _1833_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5326_ VPWR VGND _0796_ round_key[32] new_block[32] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8114_ VGND VPWR _3492_ _2632_ _2735_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8045_ VPWR VGND _3430_ block[61] round_key[61] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5257_ _0698_ _0727_ _0705_ _0626_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_4208_ VGND VPWR _3756_ _3755_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5188_ VGND VPWR _0658_ _0657_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_3_93 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_78_441 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7829_ VGND VPWR _3234_ _3232_ _3233_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_260 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4490_ VGND VPWR VPWR VGND _4018_ _4027_ _4011_ _4028_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_69_57 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_100_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6160_ _1557_ _1621_ _1389_ _1510_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5111_ VGND VPWR VGND VPWR _0562_ _0567_ _3879_ _0581_ ZI_sky130_fd_sc_hd__a21o_2
X_6091_ VPWR VGND VGND VPWR _1552_ _1553_ _1460_ ZI_sky130_fd_sc_hd__nor2_2
X_5042_ VPWR VGND VPWR VGND _0492_ _0512_ _0501_ _0491_ _0513_ ZI_sky130_fd_sc_hd__or4_2
X_6993_ VGND VPWR VPWR VGND _2443_ _2444_ _2379_ _2445_ ZI_sky130_fd_sc_hd__or3_2
X_5944_ VPWR VGND VGND VPWR _1405_ _1406_ _1404_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_47_113 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_48_614 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5875_ _1335_ _1337_ _1334_ _1336_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_4826_ VGND VPWR _0301_ _4061_ _0300_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_617 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7614_ VPWR VGND _3038_ _2732_ _0363_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7545_ VGND VPWR VPWR VGND _2973_ _2971_ _2975_ _2855_ _2974_ ZI_sky130_fd_sc_hd__o211a_2
X_4757_ VGND VPWR _0233_ _0230_ _0232_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_525 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7476_ VGND VPWR VGND VPWR _2894_ new_block[74] _2911_ _2909_ _0984_ _0053_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_70_171 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4688_ VPWR VGND VPWR VGND _0165_ _0164_ ZI_sky130_fd_sc_hd__inv_2
X_6427_ VPWR VGND _1885_ round_key[28] new_block[28] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6358_ VPWR VGND _1817_ _1816_ _1577_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_11_293 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5309_ VPWR VGND _0767_ _0779_ _0702_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_6289_ VPWR VGND VPWR VGND _1669_ _1748_ _1744_ _1458_ _1749_ ZI_sky130_fd_sc_hd__or4_2
X_8028_ VGND VPWR _3414_ _1065_ _3413_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_271 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_39_647 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_19_393 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_30_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_46_190 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_49_Left_162 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_81_458 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_39_16 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_100_490 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_58_Left_171 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_71_36 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_71_69 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5660_ VPWR VGND _1126_ round_key[52] new_block[52] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_29_157 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_84_241 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_67_Left_180 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4611_ VPWR VGND VGND VPWR _4125_ _4148_ _3872_ ZI_sky130_fd_sc_hd__nor2_2
X_5591_ VGND VPWR _1058_ _0794_ _1057_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7330_ VGND VPWR _2777_ _1146_ _2310_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4542_ VGND VPWR _4080_ _4074_ _4079_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_268 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7261_ VGND VPWR VGND VPWR _2213_ _2127_ _2302_ _2709_ ZI_sky130_fd_sc_hd__a21o_2
X_4473_ VGND VPWR VGND VPWR _4011_ _3950_ _4005_ _4010_ _3923_ _4008_ ZI_sky130_fd_sc_hd__a32o_2
X_6212_ VGND VPWR VPWR VGND _1671_ _1672_ _1670_ _1673_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_96_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7192_ VGND VPWR _2642_ _4085_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_0_485 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6143_ VPWR VGND VGND VPWR _1455_ _1604_ _1357_ ZI_sky130_fd_sc_hd__nor2_2
X_6074_ VPWR VGND VGND VPWR _1416_ _1536_ _1535_ ZI_sky130_fd_sc_hd__nor2_2
X_5025_ VPWR VGND VPWR VGND _0493_ _0495_ _0496_ _3867_ _3968_ ZI_sky130_fd_sc_hd__or4b_2
XFILLER_0_24_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_45_81 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6976_ VPWR VGND VPWR VGND _2203_ _2300_ _2202_ _2196_ _2428_ ZI_sky130_fd_sc_hd__a22o_2
X_5927_ VGND VPWR _1389_ _1388_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_35_105 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5858_ sword_ctr_reg\[1\] _1320_ sword_ctr_reg\[0\] new_block[21] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_17_Right_17 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4809_ VPWR VGND VGND VPWR _0284_ _3893_ _3939_ ZI_sky130_fd_sc_hd__nand2_2
X_5789_ VGND VPWR VGND VPWR _1252_ _0607_ _0747_ _0931_ _1251_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_90_288 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7528_ VGND VPWR _2960_ _0161_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7459_ VGND VPWR _2896_ _1888_ _2895_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_287 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_26_Right_26 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_39_411 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_27_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_41_28 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_54_414 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_54_469 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_35_661 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_41_108 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_5_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_106_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6830_ VGND VPWR VGND VPWR _2284_ _2196_ _2127_ _2132_ _2282_ _2187_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_15_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6761_ VPWR VGND _2129_ _2215_ _2163_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_8500_ VGND VPWR VPWR VGND clk _0102_ reset_n new_block[59] ZI_sky130_fd_sc_hd__dfrtp_2
X_5712_ VPWR VGND VPWR VGND _0746_ _0748_ _0592_ _0645_ _1177_ ZI_sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_53_Right_53 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6692_ VGND VPWR _2146_ _2145_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8431_ VGND VPWR VPWR VGND clk _0033_ reset_n new_block[118] ZI_sky130_fd_sc_hd__dfrtp_2
X_5643_ VGND VPWR VGND VPWR _1108_ _0582_ _0643_ _0751_ _1109_ ZI_sky130_fd_sc_hd__a31o_2
X_8362_ VGND VPWR _3716_ _2000_ _3715_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5574_ VPWR VGND VPWR VGND _0926_ _1041_ _0653_ _0833_ ZI_sky130_fd_sc_hd__or3b_2
XFILLER_0_5_599 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_53_480 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4525_ VPWR VGND _4063_ round_key[88] new_block[88] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7313_ VGND VPWR VPWR VGND _2525_ _2760_ _2070_ ZI_sky130_fd_sc_hd__and2b_2
X_8293_ VGND VPWR _3654_ _2847_ _3653_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_185 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7244_ VPWR VGND _2693_ _2692_ _2639_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_62_Right_62 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4456_ VGND VPWR VGND VPWR _3942_ _3990_ _3993_ _3992_ _3994_ ZI_sky130_fd_sc_hd__o22a_2
X_7175_ VPWR VGND _2625_ _2565_ _2311_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4387_ VGND VPWR _3925_ _3924_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_0_293 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6126_ VGND VPWR VGND VPWR _1009_ new_block[112] _1587_ _1584_ _1562_ _0027_ ZI_sky130_fd_sc_hd__o32a_2
X_6057_ VPWR VGND _1351_ _1519_ _1379_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5008_ VGND VPWR _0480_ _4066_ _4068_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_71_Right_71 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6959_ VPWR VGND _2412_ _2323_ _2310_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_48_274 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_36_469 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_106_357 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_16_182 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_80_Right_80 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_31_185 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_98_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_99_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_86_336 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_109_162 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_94_391 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_82_564 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_22_141 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_23_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5290_ VPWR VGND VPWR VGND _0743_ _0759_ _0753_ _0733_ _0760_ ZI_sky130_fd_sc_hd__or4_2
X_4310_ VPWR VGND VPWR VGND _3837_ _3847_ _3824_ _3846_ _3848_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_77_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4241_ VPWR VGND VPWR VGND _0001_ _3782_ round[1] round[0] ZI_sky130_fd_sc_hd__or3b_2
X_7931_ VPWR VGND VGND VPWR _3326_ _3324_ _3325_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_93_78 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7862_ VPWR VGND VGND VPWR _3264_ _3259_ _3263_ ZI_sky130_fd_sc_hd__nand2_2
X_7793_ VPWR VGND _3201_ _2932_ _1564_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6813_ VPWR VGND _2252_ _2267_ _2175_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_6744_ _2138_ _2198_ _2070_ _2175_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6675_ VPWR VGND VGND VPWR _3879_ _2129_ _2089_ _2094_ ZI_sky130_fd_sc_hd__nor3b_2
X_5626_ VGND VPWR VGND VPWR _0628_ _0619_ _0714_ _1090_ _1092_ _1091_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_45_277 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_91_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8414_ VGND VPWR VPWR VGND clk _0016_ reset_n new_block[101] ZI_sky130_fd_sc_hd__dfrtp_2
X_8345_ VGND VPWR _3701_ _1886_ _1894_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5557_ VPWR VGND VPWR VGND _1024_ _0610_ _0854_ ZI_sky130_fd_sc_hd__or2_2
X_8276_ VPWR VGND VPWR VGND _3575_ _3603_ _3638_ _3583_ _1891_ _3639_ ZI_sky130_fd_sc_hd__a221o_2
X_5488_ VPWR VGND VGND VPWR _0956_ _0955_ _0954_ _0953_ _0952_ _0674_ ZI_sky130_fd_sc_hd__o2111a_2
X_4508_ VPWR VGND VGND VPWR _4046_ _3794_ _3803_ ZI_sky130_fd_sc_hd__nand2_2
X_4439_ VGND VPWR VGND VPWR _3918_ _3974_ _3977_ _3976_ ZI_sky130_fd_sc_hd__a21oi_2
X_7227_ VPWR VGND VPWR VGND _2149_ _2368_ _2265_ _2300_ _2676_ ZI_sky130_fd_sc_hd__a22o_2
X_7158_ VPWR VGND VPWR VGND _2449_ _2607_ _2603_ _2474_ _2608_ ZI_sky130_fd_sc_hd__or4_2
X_7089_ VPWR VGND VPWR VGND _2282_ _2194_ _2302_ _2228_ _2540_ ZI_sky130_fd_sc_hd__a22o_2
X_6109_ VGND VPWR _1571_ _1569_ _1570_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_601 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_96_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_95_133 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_49_561 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_68_358 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_32_461 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_20_623 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_86_122 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_27_200 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4790_ VPWR VGND VPWR VGND _4031_ _4012_ _3903_ _3934_ _0265_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_7_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_55_553 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_12_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_82_361 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_12_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6460_ VGND VPWR VGND VPWR _1797_ _1521_ _1491_ _1616_ _1917_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_42_236 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6391_ VGND VPWR VGND VPWR _1427_ _1359_ _1496_ _1847_ _1849_ _1848_ ZI_sky130_fd_sc_hd__a2111o_2
X_5411_ VGND VPWR VGND VPWR _0880_ _0684_ _0582_ _0578_ _0577_ ZI_sky130_fd_sc_hd__and4_2
XFILLER_0_112_113 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5342_ VGND VPWR _0812_ _0810_ _0811_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_612 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8130_ VGND VPWR VGND VPWR _3507_ _3506_ _3505_ _3504_ ZI_sky130_fd_sc_hd__o21a_2
X_8061_ VGND VPWR _3444_ _1234_ _3443_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_177 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5273_ VGND VPWR VGND VPWR _0736_ _0735_ _0737_ _0738_ _0743_ _0742_ ZI_sky130_fd_sc_hd__a2111o_2
X_7012_ VPWR VGND VPWR VGND _2464_ _2461_ _2463_ ZI_sky130_fd_sc_hd__or2_2
X_4224_ VPWR VGND VGND VPWR _3751_ _3768_ dec_ctrl_reg\[1\] ZI_sky130_fd_sc_hd__nor2_2
X_7914_ VGND VPWR VGND VPWR _3240_ new_block[49] _3310_ _3307_ _1675_ _0092_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_78_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7845_ VPWR VGND VPWR VGND _3219_ _3159_ _3248_ _3237_ _1071_ _3249_ ZI_sky130_fd_sc_hd__a221o_2
X_4988_ VPWR VGND VPWR VGND _0459_ _3956_ _0460_ _3907_ _4037_ ZI_sky130_fd_sc_hd__or4b_2
X_7776_ VGND VPWR VPWR VGND _3184_ _1890_ _3186_ _3118_ _3185_ ZI_sky130_fd_sc_hd__o211a_2
X_6727_ VGND VPWR VGND VPWR _2181_ _2159_ _2155_ _2165_ _2180_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_61_501 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_125 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6658_ VGND VPWR _2112_ _2111_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5609_ VGND VPWR _1076_ _1060_ _1075_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_113 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_104_625 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6589_ VGND VPWR _2044_ _2042_ _2043_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8328_ VPWR VGND VPWR VGND _3521_ _3603_ _3685_ _0169_ _1575_ _3686_ ZI_sky130_fd_sc_hd__a221o_2
X_8259_ VGND VPWR _3623_ _1072_ _3622_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_21_Left_134 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_37_542 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_143 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_83_169 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_52_545 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_52_589 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_58_37 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_58_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5960_ VPWR VGND _1419_ _1422_ _1421_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5891_ VGND VPWR _1353_ _1352_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4911_ VGND VPWR _0385_ _4062_ _0141_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_155 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_59_177 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7630_ VGND VPWR VGND VPWR _3053_ _3051_ _4094_ _3052_ _2797_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_23_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4842_ VGND VPWR VGND VPWR _0317_ _0316_ _0315_ _0304_ ZI_sky130_fd_sc_hd__o21a_2
X_7561_ VGND VPWR _2989_ _2987_ _2988_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_309 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4773_ VPWR VGND VPWR VGND _0249_ round_key[66] block[66] ZI_sky130_fd_sc_hd__or2_2
XFILLER_0_55_350 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_15_225 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6512_ VGND VPWR VGND VPWR _1968_ _1546_ _1368_ _1966_ _1967_ ZI_sky130_fd_sc_hd__a211o_2
X_7492_ VGND VPWR _2926_ _1756_ _1816_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6443_ VGND VPWR _1901_ _1578_ _1690_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_11_442 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_30_239 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6374_ VPWR VGND _1833_ round_key[3] new_block[3] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5325_ VPWR VGND _0795_ round_key[37] new_block[37] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8113_ VGND VPWR VGND VPWR _3462_ new_block[3] _3491_ _3488_ _0294_ _0110_ ZI_sky130_fd_sc_hd__o32a_2
X_8044_ VPWR VGND VGND VPWR _3428_ _3429_ _0158_ ZI_sky130_fd_sc_hd__nor2_2
X_5256_ VPWR VGND VGND VPWR _0726_ _0630_ _0577_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_54_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4207_ VGND VPWR _3755_ _3754_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5187_ VPWR VGND _0599_ _0657_ _0595_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_64_80 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7828_ VPWR VGND _3233_ _2628_ _2421_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_93_445 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_81_607 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7759_ VGND VPWR _3170_ _2915_ _2898_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_96_272 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_25_501 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_37_350 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_44_309 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_4_417 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_107_260 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_64_191 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_40_515 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_107_293 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_69_36 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_0_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_40_559 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_0_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6090_ VGND VPWR _1552_ _1551_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5110_ VGND VPWR _0580_ _0579_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_85_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5041_ VPWR VGND VPWR VGND _0502_ _0511_ _0508_ _4027_ _0512_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_94_209 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6992_ VPWR VGND VPWR VGND _2177_ _2168_ _2096_ _2141_ _2444_ ZI_sky130_fd_sc_hd__a22o_2
X_5943_ VGND VPWR VPWR VGND _1319_ _1398_ _1313_ _1405_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_48_626 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5874_ _1287_ _1336_ _3755_ _1294_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_47_125 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_47_147 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7613_ VGND VPWR _3037_ _3035_ _3036_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_158 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4825_ VPWR VGND _0300_ round_key[91] new_block[91] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_90_404 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7544_ VPWR VGND VGND VPWR _2974_ _2971_ _2973_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_28_361 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4756_ VPWR VGND _0232_ _0231_ _0153_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7475_ VPWR VGND VPWR VGND _2892_ _2786_ _2910_ _2880_ _0231_ _2911_ ZI_sky130_fd_sc_hd__a221o_2
X_4687_ VGND VPWR _0164_ new_block[97] round_key[97] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6426_ VGND VPWR VPWR VGND _1884_ _1643_ _1860_ _1883_ _3756_ ZI_sky130_fd_sc_hd__o31a_2
XFILLER_0_31_537 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_70_183 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6357_ VPWR VGND _1816_ round_key[11] new_block[11] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5308_ VGND VPWR VGND VPWR _0778_ _0609_ _0600_ _0643_ _0642_ ZI_sky130_fd_sc_hd__and4_2
X_6288_ VPWR VGND VGND VPWR _1747_ _1745_ _1534_ _1491_ _1427_ _1748_ ZI_sky130_fd_sc_hd__a311o_2
X_8027_ VPWR VGND _3413_ _1068_ _0993_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5239_ VPWR VGND _0598_ _0709_ _0544_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_98_526 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_38_125 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_104_241 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_39_28 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_55_16 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_69_250 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_97_592 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_29_169 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_84_253 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_57_478 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4610_ VGND VPWR VPWR VGND _4144_ _4146_ _4139_ _4147_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_112_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5590_ VPWR VGND _1057_ round_key[35] new_block[35] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_20_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4541_ VGND VPWR _4079_ _4075_ _4078_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7260_ VGND VPWR VPWR VGND _2335_ _2707_ _2153_ _2708_ ZI_sky130_fd_sc_hd__or3_2
X_4472_ VGND VPWR _4010_ _4009_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6211_ VGND VPWR VGND VPWR _1672_ _1409_ _1368_ _1619_ _1493_ _1393_ ZI_sky130_fd_sc_hd__a32o_2
X_7191_ VPWR VGND _2641_ _2640_ _2638_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6142_ VPWR VGND VGND VPWR _1547_ _1603_ _1384_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_110_244 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6073_ VGND VPWR VPWR VGND _1393_ _1389_ _1391_ _1535_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_29_72 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5024_ VPWR VGND VGND VPWR _4110_ _3816_ _4131_ _4125_ _0495_ _0494_ ZI_sky130_fd_sc_hd__o221a_2
XFILLER_0_17_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6975_ VPWR VGND VPWR VGND _2187_ _2259_ _2174_ _2136_ _2427_ ZI_sky130_fd_sc_hd__a22o_2
X_5926_ VPWR VGND VGND VPWR _1388_ _3754_ _1348_ ZI_sky130_fd_sc_hd__nand2_2
X_5857_ VGND VPWR _1319_ _1318_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_44_651 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4808_ VGND VPWR VPWR VGND _3932_ _3887_ _0177_ _0283_ ZI_sky130_fd_sc_hd__or3_2
X_5788_ VPWR VGND VPWR VGND _0747_ _0771_ _0613_ _0702_ _1251_ ZI_sky130_fd_sc_hd__a22o_2
X_4739_ VGND VPWR VGND VPWR _3975_ _4125_ _3816_ _3916_ _0215_ ZI_sky130_fd_sc_hd__o22a_2
X_7527_ VPWR VGND _2959_ block[14] round_key[14] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7458_ VPWR VGND _2895_ _1681_ _1580_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6409_ _1308_ _1867_ _1534_ _1529_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_12_592 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7389_ VPWR VGND VPWR VGND _2797_ _2786_ _2831_ _2703_ _0367_ _2832_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_98_345 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_86_529 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_117 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_39_456 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_27_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_66_286 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_105_561 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_66_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_89_378 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_106_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6760_ VGND VPWR _2214_ _2213_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5711_ VGND VPWR VGND VPWR _1176_ _0761_ _0726_ _1175_ _0744_ ZI_sky130_fd_sc_hd__a211o_2
X_6691_ VPWR VGND VPWR VGND _2094_ _2145_ _3774_ _2089_ ZI_sky130_fd_sc_hd__or3b_2
XFILLER_0_31_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8430_ VGND VPWR VPWR VGND clk _0032_ reset_n new_block[117] ZI_sky130_fd_sc_hd__dfrtp_2
X_5642_ _0846_ _1108_ _0620_ _0654_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_13_301 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8361_ VGND VPWR _3715_ _1756_ _1899_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5573_ VPWR VGND VPWR VGND _1039_ _1040_ _1034_ _1035_ ZI_sky130_fd_sc_hd__or3b_2
X_4524_ VGND VPWR _4062_ new_block[93] round_key[93] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7312_ VGND VPWR VGND VPWR _2758_ _2187_ _2219_ _2299_ _2759_ ZI_sky130_fd_sc_hd__a31o_2
X_8292_ VGND VPWR _3653_ _2848_ _3652_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7243_ VGND VPWR _2692_ _2490_ _2691_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4455_ VGND VPWR VGND VPWR _3803_ _3857_ _3877_ _3993_ ZI_sky130_fd_sc_hd__a21o_2
X_7174_ VGND VPWR VGND VPWR _2624_ _3756_ _2623_ _2597_ ZI_sky130_fd_sc_hd__o21a_2
X_4386_ VGND VPWR VGND VPWR _3924_ _3891_ _3890_ _3885_ ZI_sky130_fd_sc_hd__and3b_2
X_6125_ VPWR VGND VPWR VGND _1281_ _0524_ _1586_ _0816_ _1585_ _1587_ ZI_sky130_fd_sc_hd__a221o_2
X_6056_ VPWR VGND VPWR VGND _1518_ _1442_ _1471_ ZI_sky130_fd_sc_hd__or2_2
XFILLER_0_56_81 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5007_ VGND VPWR _0479_ _0476_ _0478_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_337 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_72_80 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6958_ VPWR VGND _2411_ _1280_ _1198_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_48_253 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5909_ VGND VPWR _1371_ _1370_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_36_415 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6889_ VGND VPWR VGND VPWR _2341_ _2219_ _2338_ _2132_ _2342_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_76_584 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_48_297 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_91_543 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_23_109 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_32_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_86_Left_199 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_98_120 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_99_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_109_185 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_23_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_50_462 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_77_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4240_ VGND VPWR VGND VPWR _3781_ round[1] _3758_ round[0] ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_93_57 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7930_ VGND VPWR _3325_ _0242_ _3090_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7861_ VGND VPWR _3263_ _3260_ _3262_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6812_ VPWR VGND _2265_ _2266_ _2183_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_77_337 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7792_ VGND VPWR VGND VPWR _3153_ new_block[37] _3200_ _3198_ _0429_ _0080_ ZI_sky130_fd_sc_hd__o32a_2
X_6743_ VGND VPWR VGND VPWR _2197_ _2196_ _2194_ _2149_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_85_381 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6674_ VPWR VGND VGND VPWR _2128_ _3914_ _2104_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_73_532 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5625_ VPWR VGND VPWR VGND _0633_ _0787_ _0607_ _0602_ _1091_ ZI_sky130_fd_sc_hd__a22o_2
X_8413_ VGND VPWR VPWR VGND clk _0015_ reset_n new_block[100] ZI_sky130_fd_sc_hd__dfrtp_2
X_5556_ VGND VPWR VPWR VGND _1021_ _1022_ _1019_ _1023_ ZI_sky130_fd_sc_hd__or3_2
X_8344_ VGND VPWR _3700_ _3698_ _3699_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8275_ VPWR VGND _3638_ block[51] round_key[51] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5487_ VGND VPWR _0748_ _0664_ _0955_ _0666_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
XFILLER_0_41_462 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4507_ VGND VPWR VGND VPWR _4039_ _3920_ _4040_ _4043_ _4045_ _4044_ ZI_sky130_fd_sc_hd__a2111o_2
X_4438_ VGND VPWR _3976_ _3975_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7226_ VGND VPWR VGND VPWR _3776_ _2675_ _2072_ _2161_ _2089_ ZI_sky130_fd_sc_hd__and4bb_2
X_4369_ VPWR VGND VGND VPWR _3906_ _3907_ _3862_ ZI_sky130_fd_sc_hd__nor2_2
X_7157_ VGND VPWR VGND VPWR _2230_ _2107_ _2604_ _2605_ _2607_ _2606_ ZI_sky130_fd_sc_hd__a2111o_2
X_6108_ VPWR VGND _1570_ round_key[22] new_block[22] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7088_ VPWR VGND VPWR VGND _2266_ _2538_ _2261_ _2151_ _2539_ ZI_sky130_fd_sc_hd__or4_2
X_6039_ VPWR VGND VGND VPWR _1357_ _1501_ _1349_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_96_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_49_573 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_91_351 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Left_207 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_32_473 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_20_635 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_63_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_7_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_27_212 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_12_53 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6390_ VGND VPWR VGND VPWR _1848_ _1499_ _1474_ _1528_ _1523_ _1289_ ZI_sky130_fd_sc_hd__a32o_2
X_5410_ VPWR VGND VPWR VGND _0716_ _0677_ _0663_ _0570_ _0879_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_42_248 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_2_356 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5341_ VGND VPWR _0811_ new_block[62] round_key[62] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_125 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8060_ VPWR VGND _3443_ _0811_ _0801_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_100_309 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_112_169 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5272_ _0740_ _0742_ _0688_ _0741_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7011_ VGND VPWR VGND VPWR _2462_ _2118_ _2199_ _2233_ _2463_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_10_189 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4223_ VGND VPWR VGND VPWR _3748_ ready _3767_ _0004_ ZI_sky130_fd_sc_hd__a21o_2
X_7913_ VPWR VGND VPWR VGND _3309_ _3257_ _3308_ _3237_ _0911_ _3310_ ZI_sky130_fd_sc_hd__a221o_2
X_7844_ VPWR VGND _3248_ block[106] round_key[106] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_78_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7775_ VPWR VGND VGND VPWR _3185_ _1890_ _3184_ ZI_sky130_fd_sc_hd__nand2_2
X_6726_ VGND VPWR VGND VPWR _2180_ _2168_ _2150_ _2172_ _2179_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_92_137 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4987_ VPWR VGND VPWR VGND _0458_ _3923_ _4134_ _4189_ _3997_ _0459_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_46_598 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6657_ VPWR VGND VGND VPWR _2084_ _2111_ _2110_ ZI_sky130_fd_sc_hd__nor2_2
X_5608_ VGND VPWR _1075_ _1062_ _1074_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_637 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6588_ VGND VPWR _2043_ _1571_ _2003_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_473 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5539_ VGND VPWR _4103_ _4089_ _1007_ _1006_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
XFILLER_0_103_125 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8327_ VPWR VGND _3685_ block[24] round_key[24] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8258_ VGND VPWR _3622_ _0796_ _0907_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7209_ VPWR VGND VPWR VGND _2507_ _2196_ _2372_ _2327_ _2132_ _2658_ ZI_sky130_fd_sc_hd__a221o_2
X_8189_ VGND VPWR _3560_ _3085_ _3559_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_191 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_37_554 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_24_204 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_99_281 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5890_ VGND VPWR VPWR VGND _4097_ new_block[119] _1352_ _3752_ _1311_ ZI_sky130_fd_sc_hd__o211a_2
X_4910_ VGND VPWR _0384_ _0300_ _0383_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4841_ VGND VPWR VGND VPWR _0315_ _0304_ _0316_ _0158_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_87_498 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_59_189 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_28_510 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_23_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7560_ VPWR VGND _2988_ _2409_ _4087_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4772_ VPWR VGND VGND VPWR _0248_ round_key[66] block[66] ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_15_204 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6511_ VPWR VGND VPWR VGND _1332_ _1501_ _1345_ _1529_ _1967_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_43_513 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7491_ VPWR VGND _2925_ _1945_ _1885_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_15_237 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6442_ VGND VPWR _1900_ _1816_ _1899_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_365 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_3_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_23_281 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_101_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6373_ VPWR VGND _1832_ _1566_ _1564_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8112_ VPWR VGND VPWR VGND _3459_ _3490_ _3489_ _3468_ _1833_ _3491_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_2_175 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_2_197 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5324_ VPWR VGND _0794_ round_key[39] new_block[39] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8043_ VGND VPWR _3428_ _3424_ _3427_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5255_ VGND VPWR VGND VPWR _0723_ _0621_ _0725_ _0724_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_47_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4206_ VGND VPWR _3754_ _3753_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5186_ _0643_ _0656_ _0642_ _0626_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_3_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7827_ VGND VPWR _3232_ _2312_ _3231_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_435 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_65_137 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7758_ VGND VPWR VGND VPWR _3153_ new_block[34] _3169_ _3167_ _0229_ _0077_ ZI_sky130_fd_sc_hd__o32a_2
X_7689_ VGND VPWR VGND VPWR _2997_ new_block[92] _3106_ _3104_ _2624_ _0071_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_80_118 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6709_ VGND VPWR VGND VPWR _2083_ _2078_ _3850_ _2163_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_73_181 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_44_29 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_96_295 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_96_284 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_8_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_0_613 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_0_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5040_ VPWR VGND VPWR VGND _0510_ _0185_ _0509_ _4008_ _0183_ _0511_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_18_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_69 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_18_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6991_ VGND VPWR VGND VPWR _2443_ _2147_ _2138_ _2207_ _2123_ ZI_sky130_fd_sc_hd__and4_2
XFILLER_0_79_218 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5942_ VGND VPWR VPWR VGND _1393_ _1349_ _1391_ _1404_ ZI_sky130_fd_sc_hd__or3_2
X_5873_ VPWR VGND VGND VPWR _1305_ _1335_ _3879_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_75_435 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7612_ VPWR VGND _3036_ _2696_ _0489_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4824_ VGND VPWR _0299_ _0239_ _0298_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7543_ VGND VPWR _2973_ _2412_ _2972_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4755_ VPWR VGND _0231_ round_key[74] new_block[74] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_90_416 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_7_289 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_71_630 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7474_ VPWR VGND _2910_ block[10] round_key[10] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4686_ VPWR VGND _0163_ block[65] round_key[65] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6425_ VGND VPWR VGND VPWR _1882_ _1874_ _1883_ _1864_ _1658_ ZI_sky130_fd_sc_hd__nand4_2
XFILLER_0_31_549 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6356_ VGND VPWR VPWR VGND _1790_ _1814_ _1781_ _1815_ ZI_sky130_fd_sc_hd__or3_2
X_5307_ VGND VPWR VGND VPWR _0761_ _0726_ _0769_ _0773_ _0777_ _0776_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_59_81 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6287_ VGND VPWR VGND VPWR _1746_ _1444_ _1355_ _1430_ _1747_ ZI_sky130_fd_sc_hd__a31o_2
X_8026_ VGND VPWR VGND VPWR _3331_ new_block[59] _3412_ _3410_ _2545_ _0102_ ZI_sky130_fd_sc_hd__o32a_2
X_5238_ VGND VPWR VGND VPWR _0707_ _0704_ _0705_ _0706_ _0708_ ZI_sky130_fd_sc_hd__a31o_2
X_5169_ VGND VPWR _0639_ _0638_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_38_104 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_81_449 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_62_641 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_104_220 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_104_253 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_104_264 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_55_28 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_57_435 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_4_215 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_37_181 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_13_505 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4540_ VGND VPWR _4078_ _4076_ _4077_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_108_581 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_13_549 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_20_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4471_ VGND VPWR VGND VPWR _3830_ _4009_ _3844_ _3863_ _3824_ ZI_sky130_fd_sc_hd__and4bb_2
X_6210_ _1515_ _1671_ _1340_ _1474_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7190_ VGND VPWR _2640_ _1241_ _2639_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6141_ VPWR VGND VGND VPWR _1447_ _1602_ _1401_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_29_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6072_ VGND VPWR _1534_ _1424_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5023_ VGND VPWR VGND VPWR _3990_ _3988_ _3874_ _4153_ _0494_ ZI_sky130_fd_sc_hd__o22a_2
X_6974_ VPWR VGND VPWR VGND _2266_ _2159_ _2236_ _2202_ _2213_ _2426_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_0_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5925_ VPWR VGND VPWR VGND _1386_ _1381_ _1379_ _1361_ _1376_ _1387_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_48_413 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_0_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5856_ VPWR VGND VGND VPWR _3774_ _1316_ _1317_ _1318_ ZI_sky130_fd_sc_hd__nor3_2
XPHY_EDGE_ROW_3_Right_3 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4807_ VGND VPWR VGND VPWR _3918_ _3816_ _3961_ _0282_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_63_438 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5787_ VPWR VGND VPWR VGND _0761_ _1249_ _1248_ _0715_ _1250_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_16_376 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4738_ VGND VPWR VPWR VGND _0212_ _0213_ _0211_ _0214_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_44_663 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7526_ VGND VPWR VPWR VGND _2956_ _2951_ _2958_ _2855_ _2957_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_9_72 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4669_ VPWR VGND _0146_ _0145_ _4076_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7457_ VGND VPWR VGND VPWR _2894_ new_block[72] _2893_ _2890_ _0793_ _0051_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_3_281 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6408_ VGND VPWR VGND VPWR _1518_ _1397_ _1865_ _1866_ ZI_sky130_fd_sc_hd__a21o_2
X_7388_ VPWR VGND _2831_ block[35] round_key[35] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6339_ VGND VPWR VGND VPWR _1798_ _1334_ _1393_ _1389_ _1355_ _1797_ ZI_sky130_fd_sc_hd__a41o_2
X_8009_ VGND VPWR _3397_ _0806_ _1069_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_22_302 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_34_151 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_1_207 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_105_573 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_22_379 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_105_Left_218 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_89_302 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_82_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_15_97 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_18_608 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5710_ VPWR VGND VPWR VGND _0863_ _0674_ _0653_ _0675_ _0757_ _1175_ ZI_sky130_fd_sc_hd__a221o_2
X_6690_ VGND VPWR _2144_ _2143_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5641_ VGND VPWR VGND VPWR _1107_ _0747_ _0669_ _0616_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_41_600 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8360_ VGND VPWR VGND VPWR new_block[27] _3462_ _2545_ _3714_ _0134_ ZI_sky130_fd_sc_hd__o22a_2
X_5572_ VGND VPWR VPWR VGND _1036_ _0923_ _1039_ _1038_ _1037_ ZI_sky130_fd_sc_hd__o211a_2
X_8291_ VGND VPWR _3652_ _1188_ _3651_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4523_ VPWR VGND _4061_ round_key[95] new_block[95] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7311_ VGND VPWR VGND VPWR _2758_ _2222_ _2336_ _2107_ ZI_sky130_fd_sc_hd__o21a_2
X_7242_ VPWR VGND _2691_ _2011_ _1961_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_111_554 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4454_ VGND VPWR _3992_ _3991_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7173_ VPWR VGND VPWR VGND _2608_ _2622_ _2617_ _2601_ _2623_ ZI_sky130_fd_sc_hd__or4_2
X_4385_ _3803_ _3923_ _3857_ _3881_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6124_ VPWR VGND _1586_ new_block[112] round_key[112] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6055_ VPWR VGND VPWR VGND _1513_ _1516_ _1514_ _1509_ _1517_ ZI_sky130_fd_sc_hd__or4_2
X_5006_ VGND VPWR _0478_ _4073_ _0477_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6957_ VPWR VGND _2410_ _2409_ _2317_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5908_ VPWR VGND VGND VPWR _1370_ _1368_ _1369_ ZI_sky130_fd_sc_hd__nand2_2
X_6888_ VGND VPWR VGND VPWR _2340_ _2339_ _2203_ _2299_ _2341_ ZI_sky130_fd_sc_hd__a31o_2
X_5839_ VGND VPWR VGND VPWR sword_ctr_reg\[1\] sword_ctr_reg\[0\] new_block[83] _1301_
+ ZI_sky130_fd_sc_hd__nand3b_2
X_7509_ VGND VPWR _2942_ _2940_ _2941_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8489_ VGND VPWR VPWR VGND clk _0091_ reset_n new_block[48] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_31_176 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_52_29 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_67_552 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_27_449 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_109_197 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_35_482 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_105_381 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_22_187 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_26_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_93_69 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_89_132 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7860_ VGND VPWR _3262_ _2697_ _3261_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6811_ VGND VPWR _2265_ _2264_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7791_ VPWR VGND VPWR VGND _3150_ _3159_ _3199_ _3139_ _0795_ _3200_ ZI_sky130_fd_sc_hd__a221o_2
X_6742_ VGND VPWR _2196_ _2195_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6673_ VGND VPWR _2127_ _2126_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5624_ VPWR VGND VPWR VGND _0713_ _0825_ _0606_ _0731_ _1090_ ZI_sky130_fd_sc_hd__a22o_2
X_8412_ VGND VPWR VPWR VGND clk _0014_ reset_n new_block[99] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26_493 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8343_ VGND VPWR _3699_ _1575_ _1681_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5555_ VGND VPWR VPWR VGND _0727_ _0766_ _0714_ _1022_ ZI_sky130_fd_sc_hd__or3_2
X_8274_ VGND VPWR VPWR VGND _3635_ _3630_ _3637_ _3448_ _3636_ ZI_sky130_fd_sc_hd__o211a_2
X_5486_ VGND VPWR _0639_ _0727_ _0954_ _0852_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
XFILLER_0_41_474 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4506_ _3945_ _4044_ _3804_ _4010_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7225_ VGND VPWR VPWR VGND _2571_ _2673_ _2378_ _2674_ ZI_sky130_fd_sc_hd__or3_2
X_4437_ VGND VPWR VPWR VGND _3838_ _3915_ _3831_ _3975_ ZI_sky130_fd_sc_hd__or3_2
X_7156_ VGND VPWR VGND VPWR _2606_ _2132_ _2300_ _2246_ ZI_sky130_fd_sc_hd__o21a_2
X_6107_ VPWR VGND _1569_ round_key[21] new_block[21] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4368_ VGND VPWR _3906_ _3905_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_67_81 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7087_ VPWR VGND VGND VPWR _2538_ _2249_ _2328_ ZI_sky130_fd_sc_hd__nand2_2
X_4299_ VGND VPWR VPWR VGND _3835_ _3836_ _3832_ _3837_ ZI_sky130_fd_sc_hd__or3_2
X_6038_ VPWR VGND VPWR VGND _1341_ _1443_ _1346_ _1499_ _1500_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_95_113 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7989_ VGND VPWR _3379_ _1063_ _3378_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_533 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_91_363 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_32_485 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_20_658 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_63_39 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_59_349 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_94_190 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_70_503 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_70_525 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5340_ VGND VPWR _0810_ _0808_ _0809_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_137 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5271_ VPWR VGND VGND VPWR _0632_ _0741_ _0531_ ZI_sky130_fd_sc_hd__nor2_2
X_7010_ VPWR VGND VPWR VGND _2132_ _2159_ _2115_ _2155_ _2462_ ZI_sky130_fd_sc_hd__a22o_2
X_4222_ VPWR VGND VPWR VGND _3767_ dec_ctrl_reg\[1\] _3765_ dec_ctrl_reg\[0\] _3761_
+ _0002_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_37_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7912_ VGND VPWR _3309_ _3149_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_77_113 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7843_ VGND VPWR VGND VPWR _3247_ _3246_ _3245_ _3242_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_53_83 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_93_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7774_ VGND VPWR _3184_ _3181_ _3183_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4986_ VPWR VGND VPWR VGND _3911_ _3950_ _4010_ _3923_ _0458_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_46_533 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6725_ VPWR VGND _2174_ _2179_ _2178_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_6656_ VGND VPWR _2110_ _2109_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5607_ VGND VPWR _1074_ _1067_ _1073_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6587_ VGND VPWR _2042_ _1899_ _2041_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5538_ VGND VPWR _1006_ round_key[106] new_block[106] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_137 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8326_ VGND VPWR VPWR VGND _3682_ _3681_ _3684_ _0366_ _3683_ ZI_sky130_fd_sc_hd__o211a_2
X_8257_ VGND VPWR _3621_ _2848_ _3620_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7208_ VPWR VGND VPWR VGND _2651_ _2656_ _2654_ _2649_ _2657_ ZI_sky130_fd_sc_hd__or4_2
X_5469_ VGND VPWR VGND VPWR _0937_ _0729_ _0662_ _0744_ _0936_ ZI_sky130_fd_sc_hd__a211o_2
X_8188_ VGND VPWR _3559_ _0434_ _0300_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7139_ _2163_ _2589_ _2297_ _2373_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_37_500 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_96_477 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_83_105 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_24_216 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_52_514 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_52_558 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_59_113 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_90_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4840_ VGND VPWR _0315_ _0306_ _0314_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_28_522 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_28_533 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6510_ _1444_ _1966_ _1336_ _1426_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_23_97 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4771_ VGND VPWR VGND VPWR _0247_ _0246_ _0245_ _0237_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_15_216 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7490_ VGND VPWR VGND VPWR _2894_ new_block[75] _2924_ _2922_ _1054_ _0054_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_3_611 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_99_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6441_ VPWR VGND _1899_ _1898_ _1577_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_70_355 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6372_ VGND VPWR _1831_ _1563_ _1684_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5323_ VGND VPWR VPWR VGND _0760_ _0792_ _0721_ _0793_ ZI_sky130_fd_sc_hd__or3_2
X_8111_ VGND VPWR _3490_ _0161_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8042_ VGND VPWR _3427_ _3425_ _3426_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5254_ VPWR VGND VGND VPWR _0724_ _0698_ _0569_ ZI_sky130_fd_sc_hd__nand2_2
X_5185_ VGND VPWR VGND VPWR _0576_ _0593_ _0655_ _3880_ ZI_sky130_fd_sc_hd__a21oi_2
X_4205_ VGND VPWR _3753_ _3752_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7826_ VGND VPWR _3231_ _0818_ _1198_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_477 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4969_ VGND VPWR _0442_ _0439_ _0441_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7757_ VPWR VGND VPWR VGND _3150_ _3159_ _3168_ _3139_ _0985_ _3169_ ZI_sky130_fd_sc_hd__a221o_2
X_7688_ VPWR VGND VPWR VGND _2995_ _2960_ _3105_ _2984_ _0382_ _3106_ ZI_sky130_fd_sc_hd__a221o_2
X_6708_ VGND VPWR _2162_ _2129_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_34_536 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6639_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[123] sword_ctr_reg\[0\] _2093_
+ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_73_193 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_61_377 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8309_ VGND VPWR VGND VPWR _3640_ new_block[22] _3668_ _3666_ _1996_ _0129_ ZI_sky130_fd_sc_hd__o32a_2
XPHY_EDGE_ROW_110_Right_110 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_71_108 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_52_344 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_33_591 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_18_53 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6990_ VPWR VGND VGND VPWR _2124_ _2142_ _2207_ _2203_ _2282_ _2442_ ZI_sky130_fd_sc_hd__a311o_2
X_5941_ VGND VPWR VGND VPWR _1397_ _1395_ _1402_ _1403_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_34_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5872_ VPWR VGND VGND VPWR _1333_ _1334_ _3879_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_34_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_48_639 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7611_ VPWR VGND _3035_ _3034_ _2689_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4823_ VPWR VGND _0298_ _0152_ _4073_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7542_ VPWR VGND _2972_ _2691_ _2048_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4754_ VPWR VGND _0230_ round_key[79] new_block[79] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_62_108 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7473_ VGND VPWR VGND VPWR _2909_ _2908_ _2907_ _2905_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_71_642 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_71_664 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4685_ VGND VPWR _0162_ _0161_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6424_ VGND VPWR VGND VPWR _1882_ _1881_ _1878_ _1738_ _1736_ ZI_sky130_fd_sc_hd__and4_2
X_6355_ VPWR VGND VPWR VGND _1801_ _1813_ _1807_ _1799_ _1814_ ZI_sky130_fd_sc_hd__or4_2
X_6286_ VGND VPWR VGND VPWR _1487_ _1475_ _1746_ _1447_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_59_93 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5306_ VPWR VGND _0654_ _0776_ _0775_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_8025_ VPWR VGND VPWR VGND _3309_ _3367_ _3411_ _3328_ _1064_ _3412_ ZI_sky130_fd_sc_hd__a221o_2
X_5237_ VGND VPWR VGND VPWR _0707_ _0615_ _0580_ _0690_ _0666_ _0577_ ZI_sky130_fd_sc_hd__a32o_2
X_5168_ _0530_ _0638_ _3753_ _0594_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5099_ VGND VPWR _0569_ _0568_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_109_505 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_78_296 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7809_ VPWR VGND VGND VPWR _3216_ _3212_ _3215_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_46_160 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_62_664 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_18_Left_131 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_104_276 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_140 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_44_119 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_4_205 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_53_620 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_4_227 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_20_65 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4470_ VGND VPWR _4008_ _3795_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6140_ VGND VPWR VGND VPWR _1601_ _1351_ _1341_ _1546_ _1600_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_110_224 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_0_477 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6071_ VPWR VGND VPWR VGND _1532_ _1308_ _1529_ _1527_ _1499_ _1533_ ZI_sky130_fd_sc_hd__a221o_2
X_5022_ VPWR VGND VPWR VGND _0449_ _3911_ _4033_ _3926_ _4030_ _0493_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_45_40 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6973_ VPWR VGND VGND VPWR _2424_ _2423_ _2188_ _2330_ _2158_ _2425_ ZI_sky130_fd_sc_hd__a311o_2
X_5924_ VPWR VGND VGND VPWR _1385_ _1386_ _1384_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_0_53 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5855_ VPWR VGND VGND VPWR _3828_ _1317_ new_block[118] ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_0_97 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4806_ VGND VPWR VPWR VGND _0277_ _0280_ _0276_ _0281_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_90_203 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5786_ VGND VPWR VGND VPWR _0763_ _0656_ _0788_ _1249_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_9_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_43_152 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4737_ VPWR VGND VPWR VGND _4133_ _4030_ _3913_ _3926_ _0213_ ZI_sky130_fd_sc_hd__a22o_2
X_7525_ VPWR VGND VGND VPWR _2957_ _2951_ _2956_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_9_84 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_9_95 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_16_388 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4668_ VGND VPWR _0145_ _4065_ _0144_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7456_ VGND VPWR _2894_ _2799_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6407_ VGND VPWR VGND VPWR _1865_ _1522_ _1351_ _1346_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_3_293 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7387_ VGND VPWR VGND VPWR _2830_ _2829_ _2828_ _2821_ ZI_sky130_fd_sc_hd__o21a_2
X_4599_ VGND VPWR VGND VPWR _4134_ _4133_ _4136_ _4135_ ZI_sky130_fd_sc_hd__a21oi_2
X_6338_ VGND VPWR VGND VPWR _1456_ _1511_ _1401_ _1384_ _1797_ ZI_sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_101_257 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_101_268 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6269_ VPWR VGND VPWR VGND _1728_ _1521_ _1727_ _1453_ _1557_ _1729_ ZI_sky130_fd_sc_hd__a221o_2
X_8008_ VGND VPWR _3396_ _1184_ _3395_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_160 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_34_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_81_258 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_34_163 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_105_552 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_50_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_105_585 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_89_314 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_57_200 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5640_ VGND VPWR VPWR VGND _1101_ _1105_ _1099_ _1106_ ZI_sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_22_Right_22 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5571_ VPWR VGND VGND VPWR _1038_ _0616_ _0763_ ZI_sky130_fd_sc_hd__nand2_2
X_8290_ VGND VPWR _3651_ _0805_ _1126_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_174 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_53_472 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7310_ VPWR VGND VPWR VGND _2749_ _2756_ _2751_ _2747_ _2757_ ZI_sky130_fd_sc_hd__or4_2
X_4522_ VPWR VGND VPWR VGND _3964_ _4059_ _3980_ _3953_ _4060_ ZI_sky130_fd_sc_hd__or4_2
X_7241_ VGND VPWR _2690_ _2560_ _2689_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4453_ VPWR VGND VPWR VGND _3901_ _3991_ _3846_ _3837_ ZI_sky130_fd_sc_hd__or3b_2
X_7172_ VPWR VGND VGND VPWR _2621_ _2620_ _2343_ _2330_ _2214_ _2622_ ZI_sky130_fd_sc_hd__a311o_2
XFILLER_0_111_588 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4384_ VPWR VGND VGND VPWR _3921_ _3922_ _3865_ ZI_sky130_fd_sc_hd__nor2_2
X_6123_ VPWR VGND _1585_ block[16] round_key[16] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6054_ _1354_ _1516_ _1515_ _1474_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_31_Right_31 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5005_ VGND VPWR _0477_ _0149_ _0373_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_56_61 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_22_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6956_ VPWR VGND _2409_ _2011_ _1695_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_76_520 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5907_ VGND VPWR VGND VPWR _1305_ _1333_ _3796_ _1369_ ZI_sky130_fd_sc_hd__a21o_2
X_6887_ _2299_ _2340_ _2203_ _2166_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5838_ VGND VPWR VPWR VGND _1298_ _1297_ _1296_ _3822_ _1299_ _1300_ ZI_sky130_fd_sc_hd__a41oi_2
XPHY_EDGE_ROW_40_Right_40 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5769_ VGND VPWR _1233_ _0994_ _1232_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_385 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_16_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_32_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_44_483 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_44_494 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7508_ VPWR VGND _2941_ _2926_ _1898_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8488_ VGND VPWR VPWR VGND clk _0090_ reset_n new_block[47] ZI_sky130_fd_sc_hd__dfrtp_2
X_7439_ VGND VPWR _0365_ _1193_ _2878_ _2877_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
XFILLER_0_102_533 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_98_188 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_67_542 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_82_556 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_54_269 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_93_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_89_144 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_89_177 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6810_ VPWR VGND VGND VPWR _2095_ _2264_ _2117_ ZI_sky130_fd_sc_hd__nor2_2
X_7790_ VPWR VGND _3199_ block[5] round_key[5] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_9_149 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_42_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6741_ VPWR VGND _2060_ _2195_ _2139_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_42_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6672_ VPWR VGND VGND VPWR _2083_ _2126_ _3776_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_5_311 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_45_269 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8411_ VGND VPWR VPWR VGND clk _0013_ reset_n new_block[98] ZI_sky130_fd_sc_hd__dfrtp_2
X_5623_ VGND VPWR VPWR VGND _1086_ _1088_ _1085_ _1089_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_14_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8342_ VGND VPWR _3698_ _1756_ _3697_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5554_ VGND VPWR VGND VPWR _1021_ _0702_ _0675_ _0847_ _1020_ ZI_sky130_fd_sc_hd__a211o_2
X_8273_ VPWR VGND VGND VPWR _3636_ _3630_ _3635_ ZI_sky130_fd_sc_hd__nand2_2
X_5485_ VGND VPWR _0690_ _0675_ _0953_ _0651_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
X_4505_ VGND VPWR VGND VPWR _4043_ _4033_ _3945_ _4042_ _4031_ _3795_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_6_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4436_ VGND VPWR _3974_ _3973_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7224_ VPWR VGND VPWR VGND _2115_ _2154_ _2072_ _2285_ _2673_ ZI_sky130_fd_sc_hd__a22o_2
X_7155_ _2205_ _2605_ _2188_ _2208_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_4367_ VGND VPWR _3905_ _3904_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6106_ VGND VPWR _1568_ new_block[23] round_key[23] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_67_93 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7086_ VGND VPWR VPWR VGND _2534_ _2536_ _2532_ _2537_ ZI_sky130_fd_sc_hd__or3_2
X_4298_ VPWR VGND VGND VPWR _3828_ _3836_ new_block[100] ZI_sky130_fd_sc_hd__nor2_2
X_6037_ VGND VPWR _1499_ _1498_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7988_ VGND VPWR _3378_ _0800_ _0904_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_542 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_95_125 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6939_ VPWR VGND VPWR VGND _2392_ _2389_ _2391_ ZI_sky130_fd_sc_hd__or2_2
XFILLER_0_76_350 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_64_545 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_8_160 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_8_193 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_102_330 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_103_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_82_331 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_88_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5270_ VGND VPWR _0740_ _0739_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_10_136 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4221_ VPWR VGND VGND VPWR _3759_ _3767_ _3766_ ZI_sky130_fd_sc_hd__nor2_2
X_7911_ VPWR VGND _3308_ block[81] round_key[81] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7842_ VGND VPWR VGND VPWR _3245_ _3242_ _3246_ _3028_ ZI_sky130_fd_sc_hd__a21oi_2
X_4985_ VPWR VGND VPWR VGND _0454_ _0456_ _0457_ _4118_ _4152_ ZI_sky130_fd_sc_hd__or4b_2
XFILLER_0_53_95 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_93_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7773_ VGND VPWR _3183_ _1955_ _3182_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_512 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6724_ VGND VPWR _2178_ _2177_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_18_236 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_73_353 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_33_206 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_33_228 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6655_ VGND VPWR VPWR VGND _2089_ _2094_ _3774_ _2109_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_61_515 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5606_ VGND VPWR _1073_ _1070_ _1072_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6586_ VGND VPWR _2041_ _1564_ _1689_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5537_ VPWR VGND VPWR VGND _1005_ round_key[42] block[42] ZI_sky130_fd_sc_hd__or2_2
X_8325_ VPWR VGND VGND VPWR _3683_ _3681_ _3682_ ZI_sky130_fd_sc_hd__nand2_2
X_8256_ VPWR VGND _3620_ _2812_ _0911_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7207_ VPWR VGND VPWR VGND _2655_ _2599_ _2656_ _2391_ _2394_ ZI_sky130_fd_sc_hd__or4b_2
X_5468_ VGND VPWR VGND VPWR _0571_ _0754_ _0784_ _0936_ ZI_sky130_fd_sc_hd__a21o_2
X_5399_ VPWR VGND VPWR VGND _0867_ _0701_ _0765_ _0741_ _0841_ _0868_ ZI_sky130_fd_sc_hd__a221o_2
X_4419_ VGND VPWR VGND VPWR _3941_ _3905_ _3854_ _3957_ ZI_sky130_fd_sc_hd__a21o_2
X_8187_ VGND VPWR _3558_ _0148_ _3350_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7138_ _2132_ _2588_ _2126_ _2281_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7069_ VPWR VGND VPWR VGND _2517_ _2519_ _2518_ _2516_ _2520_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_69_626 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_56_309 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_52_526 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_58_29 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_87_445 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_75_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_28_545 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4770_ VGND VPWR VGND VPWR _0245_ _0237_ _0246_ _0158_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_28_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6440_ VPWR VGND _1898_ round_key[12] new_block[12] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_99_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_70_334 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6371_ VGND VPWR _1830_ _1759_ _1829_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5322_ VGND VPWR VPWR VGND _0782_ _0791_ _0777_ _0792_ ZI_sky130_fd_sc_hd__or3_2
X_8110_ VPWR VGND _3489_ block[99] round_key[99] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8041_ VGND VPWR _3426_ _0995_ _1140_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5253_ VPWR VGND VGND VPWR _0723_ _0722_ _0545_ ZI_sky130_fd_sc_hd__nand2_2
X_4204_ VPWR VGND VGND VPWR _3751_ _3752_ _3749_ ZI_sky130_fd_sc_hd__nor2_2
X_5184_ VGND VPWR _0654_ _0592_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_64_94 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7825_ VGND VPWR _3230_ _2416_ _2558_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_501 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_19_512 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7756_ VPWR VGND _3168_ block[2] round_key[2] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4968_ VPWR VGND _0441_ _0440_ _0240_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_74_640 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_34_504 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4899_ VPWR VGND _0373_ round_key[84] new_block[84] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7687_ VPWR VGND _3105_ block[92] round_key[92] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6707_ _2104_ _2161_ _3754_ _2160_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_34_548 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6638_ VGND VPWR VPWR VGND sword_ctr_reg\[0\] _2092_ new_block[59] ZI_sky130_fd_sc_hd__and2b_2
X_6569_ VGND VPWR VGND VPWR _1471_ _1522_ _1525_ _1877_ _2024_ _1969_ ZI_sky130_fd_sc_hd__a2111o_2
X_8308_ VPWR VGND VPWR VGND _3521_ _3603_ _3667_ _3583_ _1570_ _3668_ ZI_sky130_fd_sc_hd__a221o_2
X_8239_ VPWR VGND _3605_ _1061_ _0994_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_69_Right_69 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_65_651 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_110_417 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_78_Right_78 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_85_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5940_ VPWR VGND VGND VPWR _1401_ _1402_ _1399_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_87_220 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_34_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Right_87 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_87_264 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5871_ VGND VPWR VGND VPWR _1333_ _3828_ _1296_ _1297_ _1298_ _1299_ ZI_sky130_fd_sc_hd__a41o_2
X_7610_ VGND VPWR _3034_ _2547_ _3033_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_139 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4822_ VPWR VGND _0297_ _0296_ _0242_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_7_225 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7541_ VGND VPWR _2971_ _2550_ _2970_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4753_ VGND VPWR VPWR VGND _0195_ _0228_ _0190_ _0229_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_50_63 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7472_ VGND VPWR VGND VPWR _2907_ _2905_ _2908_ _2642_ ZI_sky130_fd_sc_hd__a21oi_2
X_6423_ VGND VPWR VGND VPWR _1390_ _1635_ _1482_ _1880_ _1879_ _1881_ ZI_sky130_fd_sc_hd__a2111oi_2
XFILLER_0_71_654 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_70_131 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4684_ VGND VPWR _0161_ _4092_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_96_Right_96 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_3_475 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6354_ VPWR VGND VPWR VGND _1809_ _1812_ _1810_ _1808_ _1813_ ZI_sky130_fd_sc_hd__or4_2
X_6285_ VGND VPWR VGND VPWR _1745_ _1557_ _1604_ _1491_ ZI_sky130_fd_sc_hd__o21a_2
X_5305_ VPWR VGND VGND VPWR _0775_ _0622_ _0774_ ZI_sky130_fd_sc_hd__nand2_2
X_8024_ VPWR VGND _3411_ block[59] round_key[59] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5236_ VGND VPWR _0706_ _0588_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_52_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5167_ VPWR VGND VGND VPWR _0637_ _0583_ _0626_ ZI_sky130_fd_sc_hd__nand2_2
X_5098_ VPWR VGND VGND VPWR _3774_ _0568_ _0567_ _0562_ ZI_sky130_fd_sc_hd__nor3b_2
XFILLER_0_109_517 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7808_ VGND VPWR _3215_ _3213_ _3214_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_459 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7739_ VGND VPWR _3153_ _3152_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_104_211 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_34_378 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_104_288 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_29_139 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_37_150 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_65_492 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_111_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_80_473 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_96_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_0_434 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6070_ VGND VPWR VGND VPWR _1532_ _1531_ _1444_ _1360_ _1452_ _1289_ ZI_sky130_fd_sc_hd__a32o_2
X_5021_ VGND VPWR VGND VPWR _0492_ _4110_ _3921_ _4153_ _4181_ _0188_ ZI_sky130_fd_sc_hd__o221ai_2
X_6972_ VPWR VGND VPWR VGND _2147_ _2218_ _2107_ _2204_ _2424_ ZI_sky130_fd_sc_hd__a22o_2
X_5923_ VPWR VGND VGND VPWR _1385_ _1336_ _1381_ ZI_sky130_fd_sc_hd__nand2_2
X_5854_ VGND VPWR VGND VPWR new_block[54] _3762_ _1314_ _3764_ _1316_ _1315_ ZI_sky130_fd_sc_hd__a221oi_2
X_4805_ VGND VPWR VPWR VGND _0278_ _0279_ _0176_ _0280_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_61_95 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_61_73 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5785_ VPWR VGND VPWR VGND _0739_ _0709_ _0635_ _0670_ _1248_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_90_215 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7524_ VGND VPWR _2956_ _2952_ _2955_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4736_ VPWR VGND VGND VPWR _3918_ _0212_ _3896_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_43_120 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_31_304 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_43_164 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7455_ VPWR VGND VPWR VGND _2892_ _2891_ _2857_ _2880_ _4077_ _2893_ ZI_sky130_fd_sc_hd__a221o_2
X_4667_ VPWR VGND _0144_ _0143_ _0142_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6406_ VGND VPWR VGND VPWR _1481_ _1863_ _1864_ _1342_ _1509_ ZI_sky130_fd_sc_hd__nor4_2
X_7386_ VGND VPWR VGND VPWR _2828_ _2821_ _2829_ _2642_ ZI_sky130_fd_sc_hd__a21oi_2
X_6337_ VGND VPWR VGND VPWR _1516_ _1521_ _1359_ _1427_ _1796_ ZI_sky130_fd_sc_hd__a31o_2
X_4598_ VPWR VGND VGND VPWR _4023_ _4135_ _3896_ ZI_sky130_fd_sc_hd__nor2_2
X_6268_ VPWR VGND VGND VPWR _1466_ _1728_ _1412_ ZI_sky130_fd_sc_hd__nor2_2
X_8007_ VGND VPWR _3395_ _0992_ _3394_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6199_ VPWR VGND VPWR VGND _1345_ _1528_ _1378_ _1428_ _1660_ ZI_sky130_fd_sc_hd__a22o_2
X_5219_ VPWR VGND VGND VPWR _0617_ _0689_ _0629_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_34_175 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_50_602 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_50_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_105_597 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_100_291 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_110_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5570_ VGND VPWR _0661_ _0671_ _1037_ _0859_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
XFILLER_0_31_98 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_41_613 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_41_624 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4521_ VPWR VGND VPWR VGND _4007_ _4058_ _4028_ _3996_ _4059_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_13_337 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7240_ VGND VPWR _2689_ _2309_ _2625_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4452_ VGND VPWR _3990_ _3989_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_0_253 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4383_ VPWR VGND VGND VPWR _3921_ _3894_ _3920_ ZI_sky130_fd_sc_hd__nand2_2
X_7171_ VPWR VGND VPWR VGND _2108_ _2338_ _2216_ _2229_ _2214_ _2621_ ZI_sky130_fd_sc_hd__a221o_2
X_6122_ VGND VPWR VGND VPWR _1584_ _1583_ _1582_ _1573_ ZI_sky130_fd_sc_hd__o21a_2
XPHY_EDGE_ROW_0_Left_113 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6053_ VGND VPWR _1515_ _1295_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5004_ VPWR VGND _0476_ _0308_ _4062_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_56_73 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_15_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6955_ VGND VPWR VPWR VGND _2408_ _2335_ _2351_ _2407_ _3755_ ZI_sky130_fd_sc_hd__o31a_2
X_5906_ VGND VPWR _1368_ _1367_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6886_ VGND VPWR _2339_ _2105_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5837_ VPWR VGND VGND VPWR sword_ctr_reg\[0\] sword_ctr_reg\[1\] new_block[114] _1299_
+ ZI_sky130_fd_sc_hd__nor3_2
XPHY_EDGE_ROW_46_Left_159 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5768_ VPWR VGND _1232_ _1068_ _0811_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_17_654 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8487_ VGND VPWR VPWR VGND clk _0089_ reset_n new_block[46] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7507_ VGND VPWR _2940_ _1886_ _2939_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4719_ VGND VPWR VPWR VGND _4173_ _0194_ _4007_ _0195_ ZI_sky130_fd_sc_hd__or3_2
X_7438_ VGND VPWR _2877_ _2874_ _2876_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_197 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5699_ _0615_ _1164_ _0688_ _0545_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_102_545 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7369_ VGND VPWR _2813_ _1184_ _2812_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_55_Left_168 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_105_Right_105 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_67_521 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_64_Left_177 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_22_101 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_23_613 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_2_529 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_50_421 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_112_309 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_62_281 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_77_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Left_186 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_93_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_26_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6740_ VGND VPWR _2194_ _2193_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_82_Left_195 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_42_53 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_45_237 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6671_ VGND VPWR VGND VPWR _2097_ _2073_ _2108_ _2116_ _2125_ _2124_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_42_97 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_73_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8410_ VGND VPWR VPWR VGND clk _0012_ reset_n new_block[97] ZI_sky130_fd_sc_hd__dfrtp_2
X_5622_ VGND VPWR VGND VPWR _1087_ _0704_ _0654_ _0648_ _1088_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_14_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5553_ VPWR VGND VPWR VGND _0678_ _0717_ _0615_ _0670_ _1020_ ZI_sky130_fd_sc_hd__a22o_2
X_8341_ VPWR VGND _3697_ _1759_ _1579_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_5_378 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_13_101 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_14_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4504_ VGND VPWR _4042_ _4041_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8272_ VGND VPWR _3635_ _2822_ _3634_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5484_ VGND VPWR VGND VPWR _0771_ _0859_ _0952_ _0867_ ZI_sky130_fd_sc_hd__a21oi_2
X_4435_ VGND VPWR VPWR VGND _3878_ _3929_ _3794_ _3973_ ZI_sky130_fd_sc_hd__or3_2
X_7223_ VPWR VGND VPWR VGND _2671_ _2149_ _2178_ _2187_ _2246_ _2672_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_6_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7154_ VPWR VGND _2123_ _2604_ _2236_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_4366_ VPWR VGND VPWR VGND _3901_ _3904_ _3846_ _3863_ ZI_sky130_fd_sc_hd__or3b_2
X_6105_ VGND VPWR _1567_ _1565_ _1566_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7085_ VGND VPWR VGND VPWR _2536_ _2236_ _2338_ _2303_ _2535_ ZI_sky130_fd_sc_hd__a211o_2
X_4297_ VGND VPWR VGND VPWR new_block[36] _3762_ _3833_ _3764_ _3835_ _3834_ ZI_sky130_fd_sc_hd__a221oi_2
X_6036_ _1363_ _1498_ _1312_ _1377_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_83_93 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7987_ VGND VPWR VGND VPWR _3331_ new_block[55] _3377_ _3375_ _2038_ _0098_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_49_554 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6938_ VPWR VGND VPWR VGND _2390_ _2193_ _2300_ _2285_ _2204_ _2391_ ZI_sky130_fd_sc_hd__a221o_2
X_6869_ VPWR VGND _2323_ new_block[120] round_key[120] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_64_557 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_106_169 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_103_69 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_23_498 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4220_ VPWR VGND VPWR VGND _3766_ dec_ctrl_reg\[3\] ZI_sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_90_Left_203 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7910_ VGND VPWR VPWR VGND _3305_ _3303_ _3307_ _3265_ _3306_ ZI_sky130_fd_sc_hd__o211a_2
X_7841_ VGND VPWR _3245_ _3243_ _3244_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_126 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4984_ VPWR VGND VGND VPWR _4023_ _3955_ _4181_ _3984_ _0456_ _0455_ ZI_sky130_fd_sc_hd__o221a_2
XFILLER_0_92_107 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7772_ VPWR VGND _3182_ _2000_ _1945_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6723_ VGND VPWR _2177_ _2176_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6654_ VPWR VGND _2102_ _2108_ _2107_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5605_ VGND VPWR _1072_ _0799_ _1071_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_527 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_14_410 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_26_292 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6585_ VGND VPWR _2040_ _1945_ _2039_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_82_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5536_ VPWR VGND VGND VPWR _1004_ round_key[42] block[42] ZI_sky130_fd_sc_hd__nand2_2
X_8324_ VPWR VGND _3682_ _2914_ _1832_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8255_ VGND VPWR VGND VPWR _3548_ new_block[17] _3619_ _3617_ _1675_ _0124_ ZI_sky130_fd_sc_hd__o32a_2
X_5467_ VPWR VGND VPWR VGND _0894_ _0752_ _0935_ _0772_ _0934_ ZI_sky130_fd_sc_hd__or4b_2
X_4418_ VPWR VGND VPWR VGND _3956_ _3859_ _3905_ ZI_sky130_fd_sc_hd__or2_2
X_7206_ VGND VPWR VGND VPWR _2198_ _2339_ _2572_ _2655_ ZI_sky130_fd_sc_hd__a21o_2
X_5398_ VGND VPWR VGND VPWR _0867_ _0684_ _0600_ _0582_ _0532_ ZI_sky130_fd_sc_hd__and4_2
XFILLER_0_111_183 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8186_ VGND VPWR VGND VPWR _3548_ new_block[10] _3557_ _3555_ _0984_ _0117_ ZI_sky130_fd_sc_hd__o32a_2
X_7137_ VPWR VGND VPWR VGND _2578_ _2586_ _2582_ _2577_ _2587_ ZI_sky130_fd_sc_hd__or4_2
X_4349_ VGND VPWR _3887_ _3886_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7068_ VPWR VGND VPWR VGND _2255_ _2279_ _2169_ _2281_ _2519_ ZI_sky130_fd_sc_hd__a22o_2
X_6019_ VPWR VGND VPWR VGND _1481_ _1478_ _1480_ ZI_sky130_fd_sc_hd__or2_2
XFILLER_0_9_470 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_107_445 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_45_590 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_28_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_83_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_55_332 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_99_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_70_346 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_2_112 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6370_ VGND VPWR _1829_ _1677_ _1828_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5321_ VGND VPWR VGND VPWR _0784_ _0722_ _0786_ _0789_ _0791_ _0790_ ZI_sky130_fd_sc_hd__a2111o_2
X_8040_ VGND VPWR _3425_ _0986_ _1192_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5252_ VGND VPWR _0722_ _0595_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4203_ VGND VPWR _3751_ _3750_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5183_ VPWR VGND VGND VPWR _0637_ _0653_ _0652_ ZI_sky130_fd_sc_hd__nor2_2
X_7824_ VGND VPWR VGND VPWR _3153_ new_block[40] _3229_ _3227_ _0793_ _0083_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_65_118 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4967_ VGND VPWR _0440_ _4074_ _0309_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7755_ VGND VPWR VPWR VGND _3165_ _3163_ _3167_ _3118_ _3166_ ZI_sky130_fd_sc_hd__o211a_2
X_4898_ VPWR VGND _0372_ _0371_ _0368_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7686_ VGND VPWR VGND VPWR _3104_ _3103_ _3102_ _3097_ ZI_sky130_fd_sc_hd__o21a_2
X_6706_ VGND VPWR VPWR VGND _2081_ _2080_ _2079_ _4097_ _2082_ _2160_ ZI_sky130_fd_sc_hd__a41oi_2
X_6637_ sword_ctr_reg\[1\] _2091_ sword_ctr_reg\[0\] new_block[27] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
X_6568_ VPWR VGND VPWR VGND _2016_ _2022_ _2020_ _2014_ _2023_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_6_473 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5519_ VGND VPWR _0987_ _0907_ _0986_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8307_ VPWR VGND _3667_ block[54] round_key[54] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6499_ VGND VPWR _1956_ _1564_ _1955_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8238_ VGND VPWR VGND VPWR _3548_ new_block[15] _3604_ _3601_ _1268_ _0122_ ZI_sky130_fd_sc_hd__o32a_2
X_8169_ VGND VPWR _3542_ _0297_ _3541_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_221 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_84_416 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_92_471 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_65_663 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_100_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_109_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5870_ VGND VPWR _1332_ _1331_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_34_65 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4821_ VGND VPWR _0296_ _0295_ _0148_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_87_276 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_7_204 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_68_490 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7540_ VGND VPWR _2970_ _0489_ _2308_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4752_ VPWR VGND VPWR VGND _0210_ _0227_ _0221_ _0202_ _0228_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_16_527 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_50_53 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4683_ VGND VPWR VGND VPWR _0160_ _0159_ _0157_ _0146_ ZI_sky130_fd_sc_hd__o21a_2
X_7471_ VGND VPWR _2907_ _1886_ _2906_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_121 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_3_421 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6422_ VPWR VGND VPWR VGND _1345_ _1434_ _1354_ _1438_ _1880_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_50_97 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6353_ VGND VPWR VGND VPWR _1523_ _1557_ _1482_ _1811_ _1812_ _1625_ ZI_sky130_fd_sc_hd__a2111o_2
X_6284_ VGND VPWR VGND VPWR _1744_ _1626_ _1375_ _1741_ _1743_ ZI_sky130_fd_sc_hd__a211o_2
X_5304_ VPWR VGND VGND VPWR _0774_ _0698_ _0609_ ZI_sky130_fd_sc_hd__nand2_2
X_8023_ VGND VPWR VPWR VGND _3408_ _1059_ _3410_ _3265_ _3409_ ZI_sky130_fd_sc_hd__o211a_2
X_5235_ VGND VPWR _0705_ _0600_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5166_ VPWR VGND _0633_ _0636_ _0635_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5097_ VGND VPWR VGND VPWR _3797_ _0563_ _0564_ _0565_ _0567_ _0566_ ZI_sky130_fd_sc_hd__o41ai_2
X_5999_ VPWR VGND VPWR VGND _1414_ _1461_ _1353_ _1318_ ZI_sky130_fd_sc_hd__or3b_2
XFILLER_0_109_529 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7807_ VGND VPWR _3214_ _1565_ _1895_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_81_419 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7738_ VGND VPWR _4099_ _3777_ _3152_ _3771_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
X_7669_ VGND VPWR _3088_ _3085_ _3087_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_473 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_29_118 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_57_427 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_37_162 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_111_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5020_ VPWR VGND VPWR VGND _3931_ _4150_ _4119_ _3893_ _0491_ ZI_sky130_fd_sc_hd__or4_2
X_6971_ VPWR VGND VPWR VGND _2260_ _2265_ _2123_ _2131_ _2423_ ZI_sky130_fd_sc_hd__a22o_2
X_5922_ VGND VPWR _1384_ _1383_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_29_641 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5853_ sword_ctr_reg\[1\] _1315_ sword_ctr_reg\[0\] new_block[22] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_61_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4804_ _4019_ _0279_ _3948_ _3946_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5784_ VPWR VGND VPWR VGND _0857_ _1246_ _1244_ _0679_ _1247_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_90_227 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7523_ VGND VPWR _2955_ _2953_ _2954_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4735_ _4133_ _0211_ _3891_ _3901_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_16_357 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4666_ VPWR VGND _0143_ round_key[89] new_block[89] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7454_ VGND VPWR _2892_ _2796_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7385_ VGND VPWR _2828_ _2822_ _2827_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_262 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6405_ VGND VPWR VGND VPWR _1862_ _1717_ _1863_ _1861_ ZI_sky130_fd_sc_hd__nand3_2
X_4597_ VPWR VGND VGND VPWR _3890_ _3891_ _3885_ _4134_ ZI_sky130_fd_sc_hd__nor3_2
X_6336_ VPWR VGND VPWR VGND _1421_ _1794_ _1289_ _1603_ _1795_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_12_585 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6267_ VPWR VGND VGND VPWR _1447_ _1727_ _1547_ ZI_sky130_fd_sc_hd__nor2_2
X_8006_ VGND VPWR _3394_ _0903_ _0911_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6198_ VPWR VGND VPWR VGND _1658_ _1659_ _1648_ _1651_ ZI_sky130_fd_sc_hd__or3b_2
X_5218_ VGND VPWR _0688_ _0687_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5149_ VGND VPWR _0619_ _0618_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_39_449 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_35_600 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_50_614 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_30_360 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_82_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_53_430 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_25_165 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_31_88 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4520_ VPWR VGND VPWR VGND _4045_ _4057_ _4051_ _4038_ _4058_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_103_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4451_ VGND VPWR VPWR VGND _3837_ _3915_ _3846_ _3989_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_0_221 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7170_ VPWR VGND VGND VPWR _2619_ _2349_ _2252_ _2618_ _2372_ _2620_ ZI_sky130_fd_sc_hd__a311o_2
XFILLER_0_111_524 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6121_ VGND VPWR VGND VPWR _1582_ _1573_ _1583_ _1001_ ZI_sky130_fd_sc_hd__a21oi_2
X_4382_ VPWR VGND VGND VPWR _3796_ _3920_ _3802_ _3793_ ZI_sky130_fd_sc_hd__nor3b_2
XFILLER_0_0_265 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6052_ _1358_ _1514_ _1424_ _1409_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5003_ VGND VPWR VPWR VGND _0475_ _4123_ _0465_ _0474_ _3755_ ZI_sky130_fd_sc_hd__o31a_2
XFILLER_0_56_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6954_ VPWR VGND VPWR VGND _2377_ _2406_ _2388_ _2366_ _2407_ ZI_sky130_fd_sc_hd__or4_2
X_5905_ _1347_ _1367_ _3914_ _1348_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6885_ VGND VPWR _2338_ _2136_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5836_ VPWR VGND VGND VPWR sword_ctr_reg\[0\] new_block[50] _1298_ ZI_sky130_fd_sc_hd__or2b_2
XPHY_EDGE_ROW_101_Left_214 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_63_205 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5767_ VPWR VGND _1231_ _1230_ _1229_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_17_666 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8486_ VGND VPWR VPWR VGND clk _0088_ reset_n new_block[45] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_625 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5698_ VGND VPWR VPWR VGND _1161_ _1162_ _1116_ _1163_ ZI_sky130_fd_sc_hd__or3_2
X_4718_ VPWR VGND VPWR VGND _0191_ _0193_ _0192_ _4191_ _0194_ ZI_sky130_fd_sc_hd__or4_2
X_7506_ VGND VPWR _2939_ _1569_ _1574_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7437_ VGND VPWR _2876_ _1234_ _2875_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_113 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4649_ VGND VPWR VGND VPWR _4185_ _4183_ _4186_ _4180_ _4177_ ZI_sky130_fd_sc_hd__nand4_2
X_7368_ VPWR VGND _2812_ _0912_ _0809_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_97_92 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_102_557 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6319_ VPWR VGND VGND VPWR _1778_ _1404_ _1479_ ZI_sky130_fd_sc_hd__nand2_2
X_7299_ VPWR VGND VPWR VGND _2746_ _2711_ _2713_ ZI_sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_110_Left_223 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_39_202 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_98_168 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_86_319 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_67_588 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_35_474 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_22_113 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_62_293 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_50_477 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_93_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_89_102 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_9_107 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_58_533 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_42_21 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6670_ VPWR VGND _2120_ _2124_ _2123_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5621_ VGND VPWR VGND VPWR _1087_ _0613_ _0787_ _0571_ ZI_sky130_fd_sc_hd__o21a_2
X_5552_ VPWR VGND VPWR VGND _1018_ _0953_ _1019_ _0744_ _0786_ ZI_sky130_fd_sc_hd__or4b_2
X_8340_ VGND VPWR VGND VPWR _3640_ new_block[25] _3696_ _3692_ _2408_ _0132_ ZI_sky130_fd_sc_hd__o32a_2
X_8271_ VGND VPWR _3634_ _3631_ _3633_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_113 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_14_625 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4503_ _3837_ _4041_ _3890_ _3892_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_13_146 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5483_ VPWR VGND VPWR VGND _0947_ _0950_ _0949_ _0946_ _0951_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_13_179 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4434_ VGND VPWR VGND VPWR _3969_ _3854_ _3972_ _3971_ ZI_sky130_fd_sc_hd__a21oi_2
X_7222_ VPWR VGND VPWR VGND _2285_ _2184_ _2102_ _2256_ _2671_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_1_574 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7153_ VGND VPWR VGND VPWR _2336_ _2233_ _2602_ _2381_ _2603_ _2455_ ZI_sky130_fd_sc_hd__a2111o_2
X_4365_ VGND VPWR _3903_ _3902_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6104_ VPWR VGND _1566_ round_key[0] new_block[0] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7084_ VPWR VGND VPWR VGND _2368_ _2216_ _2168_ _2208_ _2535_ ZI_sky130_fd_sc_hd__a22o_2
X_6035_ VPWR VGND VPWR VGND _1492_ _1496_ _1494_ _1488_ _1497_ ZI_sky130_fd_sc_hd__or4_2
X_4296_ sword_ctr_reg\[1\] _3834_ sword_ctr_reg\[0\] new_block[4] VPWR VGND VPWR VGND
+ ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_49_500 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_96_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7986_ VPWR VGND VPWR VGND _3309_ _3367_ _3376_ _3328_ _0993_ _3377_ ZI_sky130_fd_sc_hd__a221o_2
X_6937_ VGND VPWR VGND VPWR _2390_ _2139_ _2133_ _2105_ _2199_ ZI_sky130_fd_sc_hd__and4_2
XFILLER_0_9_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6868_ VPWR VGND _2322_ block[120] round_key[120] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5819_ VPWR VGND VPWR VGND _1281_ _0524_ _1280_ _0816_ _1279_ _1282_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_64_569 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_106_137 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6799_ VGND VPWR VGND VPWR _2253_ _2166_ _2138_ _2060_ _2252_ ZI_sky130_fd_sc_hd__and4_2
X_8469_ VGND VPWR VPWR VGND clk _0071_ reset_n new_block[92] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_477 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_103_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_55_569 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_2_305 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_11_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7840_ VGND VPWR _3244_ _2484_ _3224_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_628 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_77_105 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_53_53 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_77_138 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4983_ VGND VPWR VGND VPWR _3874_ _3978_ _3905_ _4175_ _0455_ ZI_sky130_fd_sc_hd__o22a_2
X_7771_ VGND VPWR _3181_ _1896_ _3180_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_341 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_18_216 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_92_119 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6722_ _2100_ _2176_ _2099_ _2175_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_46_558 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6653_ VGND VPWR _2107_ _2106_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_73_333 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5604_ VPWR VGND _1071_ round_key[42] new_block[42] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6584_ VPWR VGND _2039_ _1885_ _1762_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_61_539 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5535_ VGND VPWR VGND VPWR _1003_ _1002_ _1000_ _0991_ ZI_sky130_fd_sc_hd__o21a_2
X_8323_ VGND VPWR _3681_ _1950_ _3680_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8254_ VPWR VGND VPWR VGND _3575_ _3603_ _3618_ _3583_ _1759_ _3619_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_112_641 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_75_3 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5466_ VPWR VGND VPWR VGND _0718_ _0602_ _0740_ _0619_ _0706_ _0934_ ZI_sky130_fd_sc_hd__a221o_2
X_4417_ VGND VPWR _3955_ _3941_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7205_ VPWR VGND VPWR VGND _2296_ _2653_ _2652_ _2240_ _2654_ ZI_sky130_fd_sc_hd__or4_2
X_5397_ VGND VPWR VPWR VGND _0722_ _0620_ _0866_ _0654_ _0656_ ZI_sky130_fd_sc_hd__o211a_2
X_8185_ VPWR VGND VPWR VGND _3459_ _3490_ _3556_ _3468_ _1755_ _3557_ ZI_sky130_fd_sc_hd__a221o_2
X_7136_ VPWR VGND VPWR VGND _2217_ _2585_ _2584_ _2583_ _2586_ ZI_sky130_fd_sc_hd__or4_2
X_4348_ VGND VPWR VPWR VGND _3863_ _3885_ _3846_ _3886_ ZI_sky130_fd_sc_hd__or3_2
X_7067_ VGND VPWR VGND VPWR _2518_ _2193_ _2239_ _2135_ ZI_sky130_fd_sc_hd__o21a_2
X_4279_ VPWR VGND VGND VPWR _3816_ _3817_ _3795_ ZI_sky130_fd_sc_hd__nor2_2
X_6018_ VPWR VGND VGND VPWR _1479_ _1480_ _1466_ ZI_sky130_fd_sc_hd__nor2_2
X_7969_ VPWR VGND _3361_ _0373_ _0308_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_68_149 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_37_514 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_32_241 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_60_550 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_103_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_59_127 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_90_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_55_300 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_23_67 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_83_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_99_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_55_366 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_2_124 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_2_135 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5320_ _0619_ _0790_ _0577_ _0634_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_51_561 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_106_490 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5251_ VPWR VGND VPWR VGND _0681_ _0720_ _0694_ _0625_ _0721_ ZI_sky130_fd_sc_hd__or4_2
X_4202_ VPWR VGND VPWR VGND _3750_ dec_ctrl_reg\[2\] dec_ctrl_reg\[3\] ZI_sky130_fd_sc_hd__or2_2
XFILLER_0_48_53 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5182_ VPWR VGND VGND VPWR _0652_ _0532_ _0592_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_64_41 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_64_85 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7823_ VPWR VGND VPWR VGND _3219_ _3159_ _3228_ _3139_ _0903_ _3229_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_80_51 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7754_ VPWR VGND VGND VPWR _3166_ _3163_ _3165_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_46_322 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4966_ VGND VPWR _0439_ _0436_ _0438_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6705_ VGND VPWR _2159_ _2158_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_58_171 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4897_ VGND VPWR _0371_ _0369_ _0370_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7685_ VGND VPWR VGND VPWR _3102_ _3097_ _3103_ _3028_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_74_653 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_34_528 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6636_ VGND VPWR VGND VPWR _2090_ sword_ctr_reg\[0\] new_block[91] sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__and3b_2
X_6567_ VPWR VGND VPWR VGND _2021_ _1639_ _1456_ _1355_ _1346_ _2022_ ZI_sky130_fd_sc_hd__a221o_2
X_5518_ VPWR VGND _0986_ _0985_ _0794_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8306_ VGND VPWR VPWR VGND _3664_ _3659_ _3666_ _0366_ _3665_ ZI_sky130_fd_sc_hd__o211a_2
X_6498_ VGND VPWR _1955_ _1752_ _1833_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5449_ VPWR VGND VGND VPWR _0918_ round_key[41] block[41] ZI_sky130_fd_sc_hd__nand2_2
X_8237_ VPWR VGND VPWR VGND _3575_ _3603_ _3602_ _3583_ _1577_ _3604_ ZI_sky130_fd_sc_hd__a221o_2
X_8168_ VGND VPWR _3541_ _0374_ _0386_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7119_ _2127_ _2569_ _2345_ _2228_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8099_ VGND VPWR VGND VPWR _3479_ _3478_ _3477_ _3472_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_69_425 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_96_233 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_69_458 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_107_210 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_64_141 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_9_290 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_80_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_33_561 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_60_380 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_109_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4820_ VPWR VGND VPWR VGND _0295_ _4066_ ZI_sky130_fd_sc_hd__inv_2
XFILLER_0_56_631 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_7_216 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4751_ VGND VPWR VPWR VGND _0224_ _0226_ _0223_ _0227_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_7_249 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4682_ VGND VPWR VGND VPWR _0157_ _0146_ _0159_ _0158_ ZI_sky130_fd_sc_hd__a21oi_2
X_7470_ VGND VPWR _2906_ _1685_ _1752_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6421_ VPWR VGND VPWR VGND _1421_ _1511_ _1337_ _1434_ _1879_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_11_211 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6352_ VPWR VGND VGND VPWR _1552_ _1811_ _1412_ ZI_sky130_fd_sc_hd__nor2_2
X_6283_ VGND VPWR VGND VPWR _1742_ _1521_ _1523_ _1529_ _1743_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_11_255 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_11_266 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5303_ VPWR VGND VPWR VGND _0772_ _0662_ _0671_ _0757_ _0651_ _0773_ ZI_sky130_fd_sc_hd__a221o_2
X_8022_ VPWR VGND VGND VPWR _3409_ _1059_ _3408_ ZI_sky130_fd_sc_hd__nand2_2
X_5234_ VPWR VGND VGND VPWR _0704_ _0630_ _0687_ ZI_sky130_fd_sc_hd__nand2_2
X_5165_ VGND VPWR _0635_ _0634_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_38_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_75_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5096_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[111] sword_ctr_reg\[0\] _0566_
+ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_91_72 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7806_ VPWR VGND _3213_ _1569_ _1568_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5998_ VGND VPWR _1460_ _1459_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_93_225 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_59_491 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7737_ VPWR VGND VPWR VGND _3150_ _2960_ _3148_ _3139_ _0796_ _3151_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_47_664 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4949_ VGND VPWR VPWR VGND _4008_ _0421_ _0171_ _0422_ ZI_sky130_fd_sc_hd__mux2_2
X_7668_ VGND VPWR _3087_ _0311_ _3086_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6619_ VGND VPWR _2073_ _2072_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_62_645 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7599_ VGND VPWR _3024_ _2639_ _3023_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_520 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_97_520 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_53_667 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_111_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_92_291 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_21_531 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6970_ VGND VPWR VGND VPWR _1911_ new_block[121] _2422_ _2419_ _2408_ _0036_ ZI_sky130_fd_sc_hd__o32a_2
X_5921_ VGND VPWR VPWR VGND _1312_ _1363_ _1382_ _1383_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_45_98 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5852_ VPWR VGND VGND VPWR new_block[86] sword_ctr_reg\[0\] _1314_ ZI_sky130_fd_sc_hd__or2b_2
XFILLER_0_28_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4803_ VGND VPWR VGND VPWR _3992_ _4141_ _0278_ _3921_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_61_53 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5783_ VPWR VGND VPWR VGND _1245_ _0628_ _0729_ _0616_ _0651_ _1246_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_90_239 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7522_ VGND VPWR _2954_ _1565_ _1570_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4734_ VGND VPWR VGND VPWR _3931_ _0177_ _0203_ _0204_ _0210_ _0209_ ZI_sky130_fd_sc_hd__a2111o_2
X_4665_ VGND VPWR _0142_ _0141_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7453_ VPWR VGND _2891_ block[8] round_key[8] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7384_ VGND VPWR _2827_ _2824_ _2826_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_252 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6404_ VGND VPWR VGND VPWR _1609_ _1404_ _1653_ _1655_ _1424_ _1862_ ZI_sky130_fd_sc_hd__o32a_2
X_4596_ VPWR VGND VGND VPWR _3929_ _4133_ _3898_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_3_274 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6335_ VPWR VGND VGND VPWR _1794_ _1366_ _1462_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_101_92 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6266_ VGND VPWR VGND VPWR _1419_ _1359_ _1468_ _1671_ _1726_ _1725_ ZI_sky130_fd_sc_hd__a2111o_2
X_8005_ VGND VPWR VGND VPWR _3331_ new_block[57] _3393_ _3391_ _2408_ _0100_ ZI_sky130_fd_sc_hd__o32a_2
X_6197_ _1656_ _1658_ _1654_ _1657_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_5217_ VPWR VGND VGND VPWR _0687_ _3755_ _0594_ ZI_sky130_fd_sc_hd__nand2_2
X_5148_ VPWR VGND VGND VPWR _0617_ _0618_ _0531_ ZI_sky130_fd_sc_hd__nor2_2
X_5079_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] _0549_ new_block[77] ZI_sky130_fd_sc_hd__and2b_2
XFILLER_0_66_258 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_66_247 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_35_612 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_35_623 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_50_626 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_15_380 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_106_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_97_350 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_85_589 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_13_317 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_25_199 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4450_ VPWR VGND VGND VPWR _3988_ _3894_ _3959_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_53_486 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4381_ VPWR VGND VGND VPWR _3918_ _3919_ _3916_ ZI_sky130_fd_sc_hd__nor2_2
X_6120_ VPWR VGND _1582_ _1581_ _1576_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_0_277 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6051_ VGND VPWR VGND VPWR _1427_ _1346_ _1512_ _1513_ ZI_sky130_fd_sc_hd__a21o_2
X_5002_ VPWR VGND VPWR VGND _0271_ _0473_ _0470_ _3996_ _0474_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_56_97 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_88_361 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6953_ VPWR VGND VPWR VGND _2396_ _2405_ _2402_ _2392_ _2406_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_72_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5904_ VGND VPWR _1366_ _1365_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_48_203 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6884_ VGND VPWR VGND VPWR _2337_ _2336_ _2273_ _2330_ _2196_ _2252_ ZI_sky130_fd_sc_hd__a32o_2
XFILLER_0_72_85 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5835_ VGND VPWR VGND VPWR new_block[18] sword_ctr_reg\[0\] _1297_ sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__nand3_2
X_5766_ VPWR VGND _1230_ _1192_ _1058_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8485_ VGND VPWR VPWR VGND clk _0087_ reset_n new_block[44] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_155 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5697_ VPWR VGND VPWR VGND _0664_ _0701_ _0739_ _0692_ _1162_ ZI_sky130_fd_sc_hd__a22o_2
X_7505_ VGND VPWR _2938_ _1765_ _2000_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4717_ VPWR VGND VGND VPWR _3990_ _0193_ _3921_ ZI_sky130_fd_sc_hd__nor2_2
X_7436_ VGND VPWR _2875_ _0808_ _1126_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_125 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_32_637 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4648_ VPWR VGND VGND VPWR _4181_ _3918_ _4141_ _3816_ _4185_ _4184_ ZI_sky130_fd_sc_hd__o221a_2
XFILLER_0_102_503 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7367_ VPWR VGND _2811_ _0992_ _0799_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_12_361 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4579_ VGND VPWR _4116_ _3853_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_102_569 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6318_ VGND VPWR VGND VPWR _1777_ _1390_ _1606_ _1546_ ZI_sky130_fd_sc_hd__o21a_2
X_7298_ VGND VPWR VGND VPWR _4103_ new_block[126] _2745_ _2743_ _2731_ _0041_ ZI_sky130_fd_sc_hd__o32a_2
X_6249_ VPWR VGND VPWR VGND _1491_ _1639_ _1355_ _1470_ _1709_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_99_604 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_86_309 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_109_113 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_22_125 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_50_489 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_89_169 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_58_545 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_85_364 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_58_589 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5620_ VPWR VGND VPWR VGND _0650_ _0761_ _0706_ _0695_ _1086_ ZI_sky130_fd_sc_hd__a22o_2
X_5551_ VGND VPWR VGND VPWR _1018_ _0739_ _0658_ _0663_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_60_209 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8270_ VGND VPWR _3633_ _1138_ _3632_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_637 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4502_ VGND VPWR VGND VPWR _3887_ _3849_ _4040_ _3969_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_13_158 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5482_ VGND VPWR VGND VPWR _0950_ _0677_ _0545_ _0627_ _0939_ _0620_ ZI_sky130_fd_sc_hd__a32o_2
X_7221_ VPWR VGND VPWR VGND _2514_ _2669_ _2668_ _2210_ _2670_ ZI_sky130_fd_sc_hd__or4_2
X_4433_ VGND VPWR _3971_ _3970_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_1_586 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7152_ VPWR VGND _2097_ _2602_ _2231_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_4364_ _3863_ _3902_ _3846_ _3901_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7083_ VGND VPWR VGND VPWR _2534_ _2229_ _2338_ _2432_ _2533_ ZI_sky130_fd_sc_hd__a211o_2
X_6103_ VGND VPWR _1565_ _1563_ _1564_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4295_ VPWR VGND VGND VPWR new_block[68] sword_ctr_reg\[0\] _3833_ ZI_sky130_fd_sc_hd__or2b_2
X_6034_ VGND VPWR VGND VPWR _1460_ _1495_ _1496_ _1416_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_20_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_83_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7985_ VPWR VGND _3376_ block[87] round_key[87] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_96_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6936_ VGND VPWR VGND VPWR _2218_ _2203_ _2147_ _2231_ _2389_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_9_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6867_ VGND VPWR VPWR VGND _2319_ _2308_ _2321_ _1277_ _2320_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_64_515 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5818_ VGND VPWR _1281_ _4100_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_107_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6798_ VGND VPWR _2252_ _2113_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_8_185 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_51_209 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5749_ VPWR VGND VPWR VGND _1212_ _1039_ _1213_ _1207_ _1211_ ZI_sky130_fd_sc_hd__or4b_2
X_8468_ VGND VPWR VPWR VGND clk _0070_ reset_n new_block[91] ZI_sky130_fd_sc_hd__dfrtp_2
X_7419_ VGND VPWR VGND VPWR _2800_ new_block[69] _2859_ _2856_ _0429_ _0048_ ZI_sky130_fd_sc_hd__o32a_2
X_8399_ VGND VPWR VPWR VGND clk _0003_ reset_n dec_ctrl_reg\[1\] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_103_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_35_250 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_105_160 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_88_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_11_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4982_ VPWR VGND VPWR VGND _0453_ _3913_ _0218_ _4002_ _4012_ _0454_ ZI_sky130_fd_sc_hd__a221o_2
X_7770_ VGND VPWR _3180_ _1690_ _1951_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6721_ VPWR VGND VGND VPWR _3850_ _2175_ _2054_ _2059_ ZI_sky130_fd_sc_hd__nor3b_2
XFILLER_0_6_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6652_ VPWR VGND _2103_ _2106_ _2105_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_73_345 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5603_ VGND VPWR _1070_ _1068_ _1069_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_5_155 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6583_ VGND VPWR VPWR VGND _2027_ _2037_ _2023_ _2038_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_26_283 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8322_ VGND VPWR _3680_ _1580_ _1689_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_389 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5534_ VGND VPWR VGND VPWR _1000_ _0991_ _1002_ _1001_ ZI_sky130_fd_sc_hd__a21oi_2
X_8253_ VPWR VGND _3618_ block[49] round_key[49] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5465_ VGND VPWR VGND VPWR _0854_ _0630_ _0866_ _0928_ _0933_ _0932_ ZI_sky130_fd_sc_hd__a2111o_2
X_4416_ VGND VPWR _3954_ _3859_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7204_ VPWR VGND VPWR VGND _2235_ _2213_ _2167_ _2255_ _2653_ ZI_sky130_fd_sc_hd__a22o_2
X_8184_ VPWR VGND _3556_ block[74] round_key[74] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5396_ VPWR VGND _0690_ _0865_ _0695_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_7135_ VPWR VGND VPWR VGND _2302_ _2355_ _2135_ _2149_ _2585_ ZI_sky130_fd_sc_hd__a22o_2
X_4347_ VPWR VGND VPWR VGND _3883_ _3843_ _3884_ _3774_ _3885_ ZI_sky130_fd_sc_hd__or4_2
X_4278_ VPWR VGND VGND VPWR _3816_ _3804_ _3815_ ZI_sky130_fd_sc_hd__nand2_2
X_7066_ VGND VPWR VGND VPWR _2517_ _2223_ _2281_ _2204_ ZI_sky130_fd_sc_hd__o21a_2
X_6017_ VGND VPWR VPWR VGND _1393_ _1344_ _1391_ _1479_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_94_94 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7968_ VGND VPWR _3360_ _3127_ _3359_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7899_ VPWR VGND _3297_ _0147_ _4069_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6919_ VGND VPWR _2372_ _2205_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_49_386 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_91_120 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_17_250 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_91_186 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_60_573 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_103_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_87_437 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_82_120 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_83_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_36_581 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_99_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_51_573 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5250_ VGND VPWR VGND VPWR _0720_ _0703_ _0697_ _0708_ _0719_ ZI_sky130_fd_sc_hd__a211o_2
X_4201_ VPWR VGND VPWR VGND _3749_ dec_ctrl_reg\[1\] ZI_sky130_fd_sc_hd__inv_2
X_5181_ VPWR VGND VGND VPWR _0650_ _0651_ _0649_ ZI_sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_79_Left_192 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_78_415 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7822_ VPWR VGND _3228_ block[104] round_key[104] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4965_ VPWR VGND _0438_ _0437_ _0380_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_93_407 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7753_ VGND VPWR _3165_ _1757_ _3164_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6704_ VGND VPWR _2158_ _2157_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_80_63 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4896_ VGND VPWR _0370_ _4068_ _0242_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7684_ VGND VPWR _3102_ _3098_ _3101_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_27_581 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6635_ VGND VPWR VGND VPWR _3797_ _2085_ _2086_ _2087_ _2089_ _2088_ ZI_sky130_fd_sc_hd__o41ai_2
X_6566_ VGND VPWR VGND VPWR _1616_ _1308_ _1558_ _1402_ _2021_ _1432_ ZI_sky130_fd_sc_hd__a2111o_2
XFILLER_0_14_253 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8305_ VPWR VGND VGND VPWR _3665_ _3659_ _3664_ ZI_sky130_fd_sc_hd__nand2_2
X_5517_ VPWR VGND _0985_ round_key[34] new_block[34] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_42_584 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_100_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_112_461 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6497_ VGND VPWR _1954_ _1948_ _1953_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8236_ VGND VPWR _3603_ _0161_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5448_ VGND VPWR VPWR VGND _0915_ _0906_ _0917_ _0444_ _0916_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_100_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8167_ VGND VPWR VGND VPWR _3462_ new_block[8] _3540_ _3538_ _0793_ _0115_ ZI_sky130_fd_sc_hd__o32a_2
X_5379_ VPWR VGND VPWR VGND _0847_ _0628_ _0633_ _0846_ _0654_ _0848_ ZI_sky130_fd_sc_hd__a221o_2
X_8098_ VGND VPWR VGND VPWR _3477_ _3472_ _3478_ _3339_ ZI_sky130_fd_sc_hd__a21oi_2
X_7118_ _2297_ _2568_ _2339_ _2177_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7049_ VGND VPWR VGND VPWR _2499_ _2343_ _2172_ _2165_ _2500_ _2179_ ZI_sky130_fd_sc_hd__a2111o_2
XPHY_EDGE_ROW_29_Right_29 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_96_245 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_56_109 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_64_153 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_64_120 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_80_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_33_573 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_0_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_60_392 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_109_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_18_79 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4750_ VGND VPWR VPWR VGND _4039_ _0225_ _3893_ _0226_ ZI_sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_56_Right_56 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_56_654 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_55_120 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4681_ VGND VPWR _0158_ _4084_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6420_ VGND VPWR VGND VPWR _1875_ _1877_ _1878_ _1805_ _1876_ ZI_sky130_fd_sc_hd__nor4_2
XFILLER_0_43_337 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6351_ VGND VPWR VGND VPWR _1616_ _1452_ _1593_ _1637_ _1810_ _1721_ ZI_sky130_fd_sc_hd__a2111o_2
X_5302_ VPWR VGND VPWR VGND _0633_ _0771_ _0671_ _0712_ _0772_ ZI_sky130_fd_sc_hd__a22o_2
X_6282_ VGND VPWR VGND VPWR _1487_ _1538_ _1742_ _1466_ ZI_sky130_fd_sc_hd__a21oi_2
X_8021_ VGND VPWR _3408_ _3404_ _3407_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5233_ VGND VPWR VGND VPWR _0699_ _0620_ _0702_ _0703_ ZI_sky130_fd_sc_hd__a21o_2
XPHY_EDGE_ROW_87_Left_200 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_65_Right_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5164_ VPWR VGND _0557_ _0634_ _0626_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5095_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] _0565_ new_block[79] ZI_sky130_fd_sc_hd__and2b_2
XFILLER_0_91_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7805_ VGND VPWR _3212_ _2952_ _3211_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5997_ VGND VPWR VPWR VGND _1388_ _1357_ _1288_ _1459_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_93_237 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Right_74 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7736_ VGND VPWR _3150_ _3149_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_47_643 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4948_ VPWR VGND VGND VPWR _4036_ _0421_ _0182_ ZI_sky130_fd_sc_hd__nor2_2
X_4879_ VPWR VGND VPWR VGND _0351_ _0352_ _0353_ _4029_ _4054_ ZI_sky130_fd_sc_hd__or4b_2
X_7667_ VPWR VGND _3086_ _0380_ _0239_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_34_348 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6618_ VGND VPWR _2072_ _2071_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7598_ VPWR VGND _3023_ _3010_ _3022_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_42_392 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6549_ VGND VPWR _2005_ _2002_ _2004_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_83_Right_83 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8219_ VPWR VGND _3587_ _0311_ _4076_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_92_Right_92 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_53_613 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_111_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_52_167 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_21_543 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_96_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5920_ VGND VPWR VPWR VGND _1324_ _1329_ _3879_ _1382_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_0_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5851_ VGND VPWR _1313_ _1312_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_48_429 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_100_Right_100 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4802_ VGND VPWR VGND VPWR _0277_ _3946_ _4002_ _0206_ _3875_ ZI_sky130_fd_sc_hd__a211o_2
X_5782_ VGND VPWR VGND VPWR _1245_ _0717_ _0701_ _0669_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_28_175 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7521_ VGND VPWR _2953_ _1834_ _1892_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4733_ VPWR VGND VPWR VGND _0207_ _0208_ _0209_ _0205_ _0206_ ZI_sky130_fd_sc_hd__or4b_2
XFILLER_0_28_197 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7452_ VGND VPWR VGND VPWR _2890_ _2889_ _2888_ _2886_ ZI_sky130_fd_sc_hd__o21a_2
X_6403_ VGND VPWR VGND VPWR _1385_ _1366_ _1613_ _1861_ _1355_ ZI_sky130_fd_sc_hd__o2bb2a_2
X_4664_ VPWR VGND _0141_ round_key[94] new_block[94] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7383_ VGND VPWR _2826_ _2825_ _1068_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4595_ VPWR VGND VGND VPWR _4131_ _4132_ _4116_ ZI_sky130_fd_sc_hd__nor2_2
X_6334_ VGND VPWR VGND VPWR _1791_ _1529_ _1792_ _1793_ ZI_sky130_fd_sc_hd__a21o_2
X_6265_ VPWR VGND _1339_ _1725_ _1501_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_8004_ VPWR VGND VPWR VGND _3309_ _3367_ _3392_ _3328_ _0900_ _3393_ ZI_sky130_fd_sc_hd__a221o_2
X_5216_ VPWR VGND VPWR VGND _0685_ _0683_ _0677_ _0612_ _0634_ _0686_ ZI_sky130_fd_sc_hd__a221o_2
X_6196_ VGND VPWR VGND VPWR _1475_ _1405_ _1552_ _1368_ _1307_ _1657_ ZI_sky130_fd_sc_hd__o32a_2
X_5147_ VGND VPWR VPWR VGND _0537_ _0590_ _3775_ _0617_ ZI_sky130_fd_sc_hd__or3_2
X_5078_ sword_ctr_reg\[1\] _0548_ sword_ctr_reg\[0\] new_block[13] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_94_524 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_47_473 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7719_ VPWR VGND _3134_ _0230_ _0142_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_35_635 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_105_501 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_62_432 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_62_421 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_89_329 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_15_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_26_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_25_123 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_53_454 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_41_638 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4380_ VGND VPWR _3918_ _3917_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6050_ VGND VPWR VGND VPWR _1512_ _1511_ _1510_ _1491_ ZI_sky130_fd_sc_hd__o21a_2
X_5001_ VPWR VGND VPWR VGND _0471_ _0472_ _0473_ _0357_ _0424_ ZI_sky130_fd_sc_hd__or4b_2
X_6952_ VPWR VGND VPWR VGND _2291_ _2404_ _2403_ _2290_ _2405_ ZI_sky130_fd_sc_hd__or4_2
X_5903_ VGND VPWR VPWR VGND _1363_ _1364_ _1353_ _1365_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_48_215 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6883_ VGND VPWR _2336_ _2169_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_72_53 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5834_ VGND VPWR VGND VPWR sword_ctr_reg\[1\] sword_ctr_reg\[0\] new_block[82] _1296_
+ ZI_sky130_fd_sc_hd__nand3b_2
XFILLER_0_76_568 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_91_505 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5765_ VGND VPWR _1229_ _1064_ _1228_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_167 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8484_ VGND VPWR VPWR VGND clk _0086_ reset_n new_block[43] ZI_sky130_fd_sc_hd__dfrtp_2
X_5696_ VPWR VGND VPWR VGND _0683_ _0711_ _0692_ _0701_ _1161_ ZI_sky130_fd_sc_hd__a22o_2
X_4716_ VPWR VGND VGND VPWR _4114_ _0177_ _4121_ _0192_ ZI_sky130_fd_sc_hd__nor3_2
XFILLER_0_98_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7504_ VGND VPWR VGND VPWR _2894_ new_block[76] _2937_ _2935_ _1125_ _0055_ ZI_sky130_fd_sc_hd__o32a_2
X_7435_ VGND VPWR _2874_ _1228_ _2873_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_15_Left_128 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4647_ VGND VPWR VGND VPWR _3976_ _4016_ _3962_ _4023_ _4184_ ZI_sky130_fd_sc_hd__o22a_2
XFILLER_0_112_81 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_71_273 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7366_ VPWR VGND _2810_ _1135_ _1069_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_102_515 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6317_ VPWR VGND VPWR VGND _1529_ _1464_ _1337_ _1440_ _1776_ ZI_sky130_fd_sc_hd__a22o_2
X_4578_ VGND VPWR _4115_ _3978_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7297_ VPWR VGND VPWR VGND _4100_ _1959_ _2744_ _2703_ _2309_ _2745_ ZI_sky130_fd_sc_hd__a221o_2
X_6248_ VPWR VGND _1557_ _1708_ _1510_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_110_581 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6179_ VPWR VGND VPWR VGND _1501_ _1531_ _1444_ _1354_ _1640_ ZI_sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_24_Left_137 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_98_137 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_94_321 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_109_125 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_82_527 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_109_169 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_23_605 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_33_Left_146 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_22_137 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_105_364 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_30_181 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Left_155 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_26_79 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_97_181 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_58_568 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_51_Left_164 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_5_337 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5550_ VPWR VGND VPWR VGND _1012_ _1016_ _1013_ _1011_ _1017_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_5_359 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4501_ VPWR VGND VGND VPWR _3975_ _4039_ _3877_ ZI_sky130_fd_sc_hd__nor2_2
X_5481_ VGND VPWR VGND VPWR _0837_ _0621_ _0949_ _0948_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_41_435 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7220_ VGND VPWR VGND VPWR _2198_ _2128_ _2325_ _2370_ _2669_ _2431_ ZI_sky130_fd_sc_hd__a2111o_2
X_4432_ VGND VPWR VPWR VGND _3863_ _3885_ _3830_ _3970_ ZI_sky130_fd_sc_hd__or3_2
X_7151_ VGND VPWR VGND VPWR _2601_ _2159_ _2236_ _2598_ _2600_ ZI_sky130_fd_sc_hd__a211o_2
X_4363_ VGND VPWR VGND VPWR _3901_ _3843_ _3823_ _3821_ _3753_ ZI_sky130_fd_sc_hd__and4_2
XFILLER_0_1_598 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7082_ VPWR VGND VPWR VGND _2171_ _2368_ _2149_ _2259_ _2533_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_111_389 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6102_ VPWR VGND _1564_ round_key[5] new_block[5] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4294_ VGND VPWR _3832_ _3773_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_67_64 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Left_173 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6033_ VPWR VGND VGND VPWR _1495_ _1389_ _1474_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_13_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7984_ VGND VPWR VGND VPWR _3375_ _3374_ _3373_ _3370_ ZI_sky130_fd_sc_hd__o21a_2
X_6935_ VGND VPWR VGND VPWR _2378_ _2163_ _2384_ _2385_ _2388_ _2387_ ZI_sky130_fd_sc_hd__a2111o_2
X_6866_ VPWR VGND VGND VPWR _2320_ _2308_ _2319_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_76_365 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_64_527 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5817_ VPWR VGND _1280_ new_block[111] round_key[111] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_9_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6797_ VPWR VGND VPWR VGND _2250_ _2251_ _2244_ _2247_ ZI_sky130_fd_sc_hd__or3b_2
XFILLER_0_76_398 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_57_590 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5748_ VPWR VGND VPWR VGND _0943_ _0930_ _0946_ _0853_ _1212_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_106_106 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_106_117 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_107_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8536_ VGND VPWR VPWR VGND clk _0138_ reset_n new_block[31] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_72_571 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5679_ VPWR VGND _1145_ block[44] round_key[44] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_102_301 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8467_ VGND VPWR VPWR VGND clk _0069_ reset_n new_block[90] ZI_sky130_fd_sc_hd__dfrtp_2
X_7418_ VPWR VGND VPWR VGND _2797_ _2858_ _2857_ _2703_ _4068_ _2859_ ZI_sky130_fd_sc_hd__a221o_2
X_8398_ VPWR VGND VPWR VGND dec_ctrl_reg\[0\] reset_n _0002_ clk ZI_sky130_fd_sc_hd__dfstp_2
X_7349_ VPWR VGND _2795_ block[32] round_key[32] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_95_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_55_505 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_103_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_23_424 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_35_262 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_112_109 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_10_118 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_53_33 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4981_ VPWR VGND VGND VPWR _3982_ _0453_ _3859_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_98_490 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_6720_ VGND VPWR _2174_ _2173_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6651_ _2104_ _2105_ _3753_ _2083_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_6_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5602_ VPWR VGND _1069_ _0900_ _0811_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6582_ VPWR VGND VPWR VGND _2029_ _2036_ _2033_ _1933_ _2037_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_6_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5533_ VGND VPWR _1001_ _4085_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_14_402 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8321_ VGND VPWR VGND VPWR _3640_ new_block[23] _3679_ _3675_ _2038_ _0130_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_41_210 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_103_109 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8252_ VGND VPWR VPWR VGND _3615_ _3614_ _3617_ _3448_ _3616_ ZI_sky130_fd_sc_hd__o211a_2
X_5464_ VPWR VGND VGND VPWR _0931_ _0930_ _0654_ _0722_ _0648_ _0932_ ZI_sky130_fd_sc_hd__a311o_2
XFILLER_0_111_120 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_78_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5395_ VPWR VGND VPWR VGND _0607_ _0671_ _0658_ _0669_ _0864_ ZI_sky130_fd_sc_hd__a22o_2
X_8183_ VGND VPWR VGND VPWR _3555_ _3554_ _3553_ _3550_ ZI_sky130_fd_sc_hd__o21a_2
X_7203_ VPWR VGND VPWR VGND _2435_ _2123_ _2148_ _2111_ _2141_ _2652_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_78_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4415_ VPWR VGND VPWR VGND _3937_ _3952_ _3944_ _3909_ _3953_ ZI_sky130_fd_sc_hd__or4_2
X_7134_ VPWR VGND VPWR VGND _2223_ _2184_ _2072_ _2143_ _2584_ ZI_sky130_fd_sc_hd__a22o_2
X_4346_ VPWR VGND VGND VPWR _3828_ _3884_ new_block[103] ZI_sky130_fd_sc_hd__nor2_2
X_7065_ VPWR VGND VPWR VGND _2183_ _2201_ _2123_ _2143_ _2516_ ZI_sky130_fd_sc_hd__a22o_2
X_4277_ VPWR VGND VGND VPWR _3796_ _3809_ _3814_ _3815_ ZI_sky130_fd_sc_hd__nor3_2
X_6016_ VPWR VGND VGND VPWR _1473_ _1478_ _1401_ ZI_sky130_fd_sc_hd__nor2_2
X_7967_ VGND VPWR _3359_ _0150_ _0431_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_37_505 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6918_ VPWR VGND VPWR VGND _2371_ _2369_ _2370_ ZI_sky130_fd_sc_hd__or2_2
X_7898_ VGND VPWR _3296_ _4064_ _3295_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_462 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6849_ VGND VPWR VGND VPWR _2097_ _2285_ _2302_ _2213_ _2303_ ZI_sky130_fd_sc_hd__o22a_2
XFILLER_0_92_622 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_91_154 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_91_132 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_17_262 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_91_165 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8519_ VGND VPWR VPWR VGND clk _0121_ reset_n new_block[14] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_91_198 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_107_Left_220 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_103_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_2_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_102_186 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_102_197 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_87_449 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_67_151 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_82_132 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_51_541 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4200_ VPWR VGND VPWR VGND _0000_ _3748_ ZI_sky130_fd_sc_hd__inv_2
X_5180_ VGND VPWR VPWR VGND _0530_ _0576_ _3775_ _0650_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_48_99 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_3_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7821_ VGND VPWR VPWR VGND _3225_ _3222_ _3227_ _3118_ _3226_ ZI_sky130_fd_sc_hd__o211a_2
X_4964_ VGND VPWR _0437_ _4062_ _0382_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7752_ VGND VPWR _3164_ _1681_ _1764_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_75 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6703_ VGND VPWR _2157_ _2156_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4895_ VPWR VGND _0369_ _0306_ _4067_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7683_ VGND VPWR _3101_ _3099_ _3100_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_97 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6634_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[122] sword_ctr_reg\[0\] _2088_
+ ZI_sky130_fd_sc_hd__or3_2
X_6565_ VGND VPWR VGND VPWR _2020_ _1440_ _1453_ _2017_ _2019_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_89_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8304_ VGND VPWR _3664_ _3661_ _3663_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_265 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6496_ VGND VPWR _1953_ _1950_ _1952_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5516_ VGND VPWR VPWR VGND _0938_ _0983_ _0933_ _0984_ ZI_sky130_fd_sc_hd__or3_2
X_5447_ VPWR VGND VGND VPWR _0916_ _0906_ _0915_ ZI_sky130_fd_sc_hd__nand2_2
X_8235_ VPWR VGND _3602_ block[79] round_key[79] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_100_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_112_473 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_100_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8166_ VPWR VGND VPWR VGND _3459_ _3490_ _3539_ _3468_ _1579_ _3540_ ZI_sky130_fd_sc_hd__a221o_2
X_5378_ _0785_ _0847_ _0754_ _0722_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8097_ VGND VPWR _3477_ _3473_ _3476_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7117_ VGND VPWR VGND VPWR _2567_ _2202_ _2213_ _2302_ ZI_sky130_fd_sc_hd__o21a_2
X_4329_ VGND VPWR VGND VPWR _3867_ _3845_ _3817_ _3855_ _3866_ ZI_sky130_fd_sc_hd__a211o_2
X_7048_ VPWR VGND VPWR VGND _2159_ _2330_ _2150_ _2132_ _2499_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_49_162 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_49_184 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_100_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_103_495 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_109_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_56_600 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_56_666 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_55_143 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_43_316 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4680_ VGND VPWR _0157_ _0151_ _0156_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_165 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_36_390 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6350_ VPWR VGND VPWR VGND _1809_ _1502_ _1512_ ZI_sky130_fd_sc_hd__or2_2
X_5301_ VGND VPWR _0771_ _0770_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6281_ _1438_ _1741_ _1424_ _1434_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8020_ VGND VPWR _3407_ _2810_ _3406_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5232_ VGND VPWR _0702_ _0701_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5163_ VPWR VGND VGND VPWR _0632_ _0633_ _0630_ ZI_sky130_fd_sc_hd__nor2_2
X_5094_ sword_ctr_reg\[1\] _0564_ sword_ctr_reg\[0\] new_block[15] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
X_7804_ VGND VPWR _3211_ _1899_ _1945_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5996_ VGND VPWR VGND VPWR _1458_ _1452_ _1440_ _1454_ _1457_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_93_216 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_93_249 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7735_ VGND VPWR VGND VPWR _3149_ _4099_ _3771_ _3777_ ZI_sky130_fd_sc_hd__o21a_2
X_4947_ VPWR VGND VPWR VGND _4111_ _0419_ _4143_ _3943_ _0420_ ZI_sky130_fd_sc_hd__or4_2
X_4878_ VPWR VGND VGND VPWR _3999_ _3984_ _3982_ _3974_ _0352_ _3957_ ZI_sky130_fd_sc_hd__o221a_2
X_7666_ VGND VPWR _3085_ _0155_ _3084_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6617_ VPWR VGND _2060_ _2071_ _2070_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_61_113 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7597_ VGND VPWR _3022_ _1146_ _2315_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_146 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6548_ VPWR VGND _2004_ _2003_ _1563_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6479_ VPWR VGND VPWR VGND _1410_ _1935_ _1934_ _1406_ _1936_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_30_533 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_30_599 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8218_ VPWR VGND _3586_ _0514_ _3345_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8149_ VGND VPWR _3524_ _2734_ _3523_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_69_268 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_84_249 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_20_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_111_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_29_57 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5850_ VGND VPWR VGND VPWR _1312_ _1311_ _4097_ new_block[119] _3752_ ZI_sky130_fd_sc_hd__o211ai_2
XFILLER_0_75_205 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_0_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_29_655 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4801_ VPWR VGND VPWR VGND _0275_ _4042_ _0218_ _4134_ _3926_ _0276_ ZI_sky130_fd_sc_hd__a221o_2
X_5781_ VPWR VGND VPWR VGND _1243_ _0706_ _0763_ _0661_ _0731_ _1244_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_16_305 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_28_154 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7520_ VGND VPWR _2952_ _1680_ _2039_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4732_ VGND VPWR VPWR VGND _3849_ _3939_ _3930_ _0208_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_28_187 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_43_102 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7451_ VGND VPWR VGND VPWR _2888_ _2886_ _2889_ _2642_ ZI_sky130_fd_sc_hd__a21oi_2
X_4663_ VGND VPWR VPWR VGND _0140_ _4123_ _4157_ _0139_ _3756_ ZI_sky130_fd_sc_hd__o31a_2
X_6402_ VPWR VGND VPWR VGND _1850_ _1859_ _1852_ _1846_ _1860_ ZI_sky130_fd_sc_hd__or4_2
X_7382_ VGND VPWR _2825_ _0809_ _0993_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_360 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4594_ VGND VPWR _4131_ _4036_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_71_488 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6333_ VGND VPWR VGND VPWR _1792_ _1639_ _1501_ _1470_ ZI_sky130_fd_sc_hd__o21a_2
X_6264_ VPWR VGND VPWR VGND _1706_ _1723_ _1711_ _1703_ _1724_ ZI_sky130_fd_sc_hd__or4_2
X_8003_ VPWR VGND _3392_ block[57] round_key[57] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5215_ VGND VPWR VGND VPWR _0685_ _0569_ _0595_ _0684_ _0591_ ZI_sky130_fd_sc_hd__and4_2
XFILLER_0_86_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6195_ VGND VPWR VGND VPWR _1466_ _1655_ _1419_ _1656_ _1351_ ZI_sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_43_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5146_ VGND VPWR _0616_ _0615_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5077_ VGND VPWR VGND VPWR _0547_ new_block[45] sword_ctr_reg\[1\] sword_ctr_reg\[0\]
+ ZI_sky130_fd_sc_hd__and3b_2
XFILLER_0_66_205 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5979_ _1333_ _1441_ _3914_ _1392_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_109_307 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_66_238 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7718_ VGND VPWR _3133_ _4066_ _0431_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7649_ VGND VPWR VPWR VGND _3068_ _3066_ _3070_ _2855_ _3069_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_62_477 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_50_639 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_42_190 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_15_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_57_238 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_26_625 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_25_135 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_108_373 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_53_499 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_111_505 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5000_ VPWR VGND VGND VPWR _4050_ _4160_ _4193_ _0282_ _0472_ ZI_sky130_fd_sc_hd__and4b_2
X_6951_ VGND VPWR VGND VPWR _2404_ _2281_ _2162_ _2256_ _2260_ _2207_ ZI_sky130_fd_sc_hd__a32o_2
X_5902_ VPWR VGND VPWR VGND _1329_ _1364_ _3879_ _1324_ ZI_sky130_fd_sc_hd__or3b_2
XFILLER_0_48_227 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6882_ VPWR VGND VGND VPWR _2329_ _2332_ _2334_ _2335_ ZI_sky130_fd_sc_hd__nor3_2
X_5833_ VPWR VGND VGND VPWR _1294_ _1295_ _3787_ ZI_sky130_fd_sc_hd__nor2_2
X_5764_ VPWR VGND _1228_ _1137_ _0902_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7503_ VPWR VGND VPWR VGND _2892_ _2786_ _2936_ _2880_ _0376_ _2937_ ZI_sky130_fd_sc_hd__a221o_2
X_8483_ VGND VPWR VPWR VGND clk _0085_ reset_n new_block[42] ZI_sky130_fd_sc_hd__dfrtp_2
X_4715_ VPWR VGND VGND VPWR _3882_ _0191_ _3872_ ZI_sky130_fd_sc_hd__nor2_2
X_5695_ VPWR VGND VPWR VGND _1159_ _0846_ _0710_ _0757_ _0717_ _1160_ ZI_sky130_fd_sc_hd__a221o_2
X_7434_ VGND VPWR _2873_ _0811_ _0993_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4646_ VPWR VGND VGND VPWR _3998_ _3816_ _4025_ _3872_ _4183_ _4182_ ZI_sky130_fd_sc_hd__o221a_2
XFILLER_0_4_585 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_31_138 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4577_ VGND VPWR _4114_ _3865_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_102_527 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7365_ VGND VPWR VGND VPWR _2800_ new_block[65] _2809_ _2807_ _0140_ _0044_ ZI_sky130_fd_sc_hd__o32a_2
X_6316_ VPWR VGND VPWR VGND _1773_ _1774_ _1626_ _1534_ _1775_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_97_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7296_ VPWR VGND _2744_ block[126] round_key[126] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6247_ VPWR VGND VGND VPWR _1460_ _1707_ _1609_ ZI_sky130_fd_sc_hd__nor2_2
X_6178_ VGND VPWR _1639_ _1489_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5129_ _0537_ _0599_ _3752_ _0590_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_99_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_54_208 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_23_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_50_414 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_30_193 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_97_193 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_85_333 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_42_68 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5480_ VPWR VGND VPWR VGND _0643_ _0887_ _0948_ _0886_ _0642_ ZI_sky130_fd_sc_hd__or4b_2
X_4500_ VPWR VGND VPWR VGND _4032_ _4037_ _4034_ _4029_ _4038_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_13_127 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4431_ VGND VPWR _3969_ _3942_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_101_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4362_ VPWR VGND VGND VPWR _3860_ _3900_ _3878_ ZI_sky130_fd_sc_hd__nor2_2
X_7150_ VGND VPWR VGND VPWR _2599_ _2150_ _2600_ _2149_ ZI_sky130_fd_sc_hd__a21bo_2
XFILLER_0_67_32 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7081_ VPWR VGND VPWR VGND _2531_ _2259_ _2171_ _2372_ _2230_ _2532_ ZI_sky130_fd_sc_hd__a221o_2
X_6101_ VGND VPWR _1563_ new_block[6] round_key[6] VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4293_ VGND VPWR _3831_ _3830_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6032_ VGND VPWR VGND VPWR _1494_ _1493_ _1470_ _1350_ ZI_sky130_fd_sc_hd__o21a_2
X_7983_ VGND VPWR VGND VPWR _3373_ _3370_ _3374_ _3339_ ZI_sky130_fd_sc_hd__a21oi_2
X_6934_ VGND VPWR VGND VPWR _2386_ _2219_ _2372_ _2159_ _2387_ ZI_sky130_fd_sc_hd__a31o_2
X_6865_ VGND VPWR _2319_ _2314_ _2318_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5816_ VPWR VGND _1279_ block[47] round_key[47] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6796_ VGND VPWR VGND VPWR _2250_ _2249_ _2248_ _2225_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_76_388 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_44_230 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_106_129 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8535_ VGND VPWR VPWR VGND clk _0137_ reset_n new_block[30] ZI_sky130_fd_sc_hd__dfrtp_2
X_5747_ VGND VPWR VGND VPWR _1210_ _1208_ _1211_ _0923_ ZI_sky130_fd_sc_hd__a21oi_2
X_8466_ VGND VPWR VPWR VGND clk _0068_ reset_n new_block[89] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_72_583 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5678_ VGND VPWR VGND VPWR _1144_ _1143_ _1142_ _1130_ ZI_sky130_fd_sc_hd__o21a_2
X_7417_ VPWR VGND _2858_ block[37] round_key[37] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4629_ VGND VPWR VGND VPWR _3933_ _4021_ _3954_ _4141_ _4166_ ZI_sky130_fd_sc_hd__o22a_2
X_8397_ VGND VPWR VGND VPWR _3461_ new_block[31] _3747_ _3745_ _2775_ _0138_ ZI_sky130_fd_sc_hd__o32a_2
X_7348_ VGND VPWR VPWR VGND _2792_ _2789_ _2794_ _1277_ _2793_ ZI_sky130_fd_sc_hd__o211a_2
X_7279_ VGND VPWR VGND VPWR _2727_ _2222_ _2171_ _2174_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_95_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_55_517 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_63_561 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_50_233 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_105_195 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_37_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_37_79 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_53_45 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4980_ VPWR VGND VPWR VGND _0451_ _4155_ _0452_ _0184_ _0450_ ZI_sky130_fd_sc_hd__or4b_2
X_6650_ VGND VPWR VPWR VGND _2076_ _2075_ _2074_ _3828_ _2077_ _2104_ ZI_sky130_fd_sc_hd__a41oi_2
XFILLER_0_73_303 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_6_625 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6581_ VGND VPWR VGND VPWR _2036_ _1428_ _1440_ _1621_ _2035_ ZI_sky130_fd_sc_hd__a211o_2
X_5601_ VPWR VGND _1068_ round_key[51] new_block[51] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5532_ VGND VPWR _1000_ _0995_ _0999_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8320_ VPWR VGND VGND VPWR _3678_ _3458_ _0162_ _3676_ _3677_ _3679_ ZI_sky130_fd_sc_hd__a311o_2
X_8251_ VPWR VGND VGND VPWR _3616_ _3614_ _3615_ ZI_sky130_fd_sc_hd__nand2_2
X_5463_ VPWR VGND VGND VPWR _0724_ _0931_ _0652_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_10_620 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5394_ VPWR VGND _0746_ _0863_ _0627_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_4414_ VGND VPWR VGND VPWR _3952_ _3898_ _3951_ _3947_ ZI_sky130_fd_sc_hd__o21a_2
X_7202_ VGND VPWR VGND VPWR _2650_ _2343_ _2229_ _2214_ _2651_ ZI_sky130_fd_sc_hd__a31o_2
X_8182_ VGND VPWR VGND VPWR _3553_ _3550_ _3554_ _3339_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_111_132 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_78_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_111_165 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7133_ VPWR VGND _2227_ _2583_ _2208_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_78_97 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4345_ VPWR VGND VPWR VGND _3818_ _3764_ _3883_ _3819_ _3820_ ZI_sky130_fd_sc_hd__a211oi_2
X_7064_ VPWR VGND VPWR VGND _2509_ _2514_ _2511_ _2506_ _2515_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_94_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4276_ VGND VPWR VGND VPWR _3788_ _3810_ _3811_ _3812_ _3814_ _3813_ ZI_sky130_fd_sc_hd__o41ai_2
X_6015_ VPWR VGND VPWR VGND _1476_ _1332_ _1471_ _1355_ _1470_ _1477_ ZI_sky130_fd_sc_hd__a221o_2
X_7966_ VGND VPWR _3358_ _0312_ _0435_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6917_ VGND VPWR VGND VPWR _2370_ _2255_ _2279_ _2223_ ZI_sky130_fd_sc_hd__o21a_2
X_7897_ VGND VPWR _3295_ _4073_ _0150_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_76_141 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6848_ VGND VPWR _2302_ _2141_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_64_325 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_92_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_91_144 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_17_274 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_45_561 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6779_ VGND VPWR _2233_ _2115_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8518_ VGND VPWR VPWR VGND clk _0120_ reset_n new_block[13] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_266 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8449_ VGND VPWR VPWR VGND clk _0051_ reset_n new_block[72] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_99_255 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_99_299 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_23_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_95_494 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_3_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_82_188 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_23_277 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_51_586 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_48_67 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7820_ VPWR VGND VGND VPWR _3226_ _3222_ _3225_ ZI_sky130_fd_sc_hd__nand2_2
X_4963_ VPWR VGND _0436_ _0435_ _0434_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7751_ VGND VPWR _3163_ _3161_ _3162_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7682_ VPWR VGND _3100_ _0386_ _0376_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6702_ _2100_ _2156_ _2099_ _2133_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6633_ VGND VPWR VPWR VGND sword_ctr_reg\[0\] _2087_ new_block[58] ZI_sky130_fd_sc_hd__and2b_2
X_4894_ VGND VPWR _0368_ _4066_ _0367_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_645 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_73_144 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_27_561 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6564_ VGND VPWR VGND VPWR _2018_ _1344_ _1522_ _1381_ _2019_ ZI_sky130_fd_sc_hd__a31o_2
X_8303_ VGND VPWR _3663_ _1182_ _3662_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6495_ VGND VPWR _1952_ _1763_ _1951_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5515_ VPWR VGND VPWR VGND _0962_ _0982_ _0969_ _0957_ _0983_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_14_277 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5446_ VPWR VGND _0915_ _0914_ _0910_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_8234_ VGND VPWR VPWR VGND _3599_ _3596_ _3601_ _3448_ _3600_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_100_625 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5377_ VGND VPWR _0846_ _0785_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8165_ VPWR VGND _3539_ block[72] round_key[72] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7116_ VGND VPWR VGND VPWR _1911_ new_block[123] _2566_ _2563_ _2545_ _0038_ ZI_sky130_fd_sc_hd__o32a_2
X_8096_ VGND VPWR _3476_ _3474_ _3475_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4328_ VGND VPWR VGND VPWR _3862_ _3859_ _3866_ _3865_ ZI_sky130_fd_sc_hd__a21oi_2
X_7047_ VGND VPWR VGND VPWR _1911_ new_block[122] _2498_ _2495_ _2483_ _0037_ ZI_sky130_fd_sc_hd__o32a_2
X_4259_ VGND VPWR _3797_ _3788_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7949_ VPWR VGND VPWR VGND _3309_ _3257_ _3342_ _3328_ _1126_ _3343_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_107_202 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_64_111 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_107_235 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_92_486 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_80_626 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_33_520 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_20_203 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_18_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_109_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_75_409 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_56_612 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_51_350 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5300_ _0643_ _0770_ _0642_ _0568_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_6280_ VPWR VGND VPWR VGND _1730_ _1739_ _1732_ _1726_ _1740_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_11_225 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_59_44 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5231_ VGND VPWR _0701_ _0700_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5162_ VGND VPWR _0632_ _0631_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5093_ VGND VPWR VGND VPWR _0563_ new_block[47] sword_ctr_reg\[1\] sword_ctr_reg\[0\]
+ ZI_sky130_fd_sc_hd__and3b_2
XFILLER_0_75_87 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_75_65 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7803_ VGND VPWR VGND VPWR _3153_ new_block[38] _3210_ _3208_ _0475_ _0081_ ZI_sky130_fd_sc_hd__o32a_2
X_5995_ VGND VPWR VGND VPWR _1457_ _1438_ _1289_ _1456_ _1427_ _1340_ ZI_sky130_fd_sc_hd__a32o_2
X_7734_ VPWR VGND _3148_ block[0] round_key[0] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4946_ VPWR VGND VPWR VGND _4013_ _3925_ _3903_ _3923_ _0419_ ZI_sky130_fd_sc_hd__a22o_2
X_7665_ VPWR VGND _3084_ _0230_ _4078_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4877_ VGND VPWR VGND VPWR _3910_ _3931_ _0350_ _4190_ _0351_ _0207_ ZI_sky130_fd_sc_hd__a2111o_2
X_7596_ VGND VPWR _3021_ _2626_ _3020_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6616_ VPWR VGND VPWR VGND _2064_ _2063_ _2070_ _3787_ _2069_ ZI_sky130_fd_sc_hd__a211oi_2
XFILLER_0_6_296 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6547_ VGND VPWR _2003_ _1683_ _1895_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_169 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_30_545 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6478_ VPWR VGND VPWR VGND _1345_ _1409_ _1359_ _1499_ _1935_ ZI_sky130_fd_sc_hd__a22o_2
X_8217_ VGND VPWR VGND VPWR _3548_ new_block[13] _3585_ _3582_ _1181_ _0120_ ZI_sky130_fd_sc_hd__o32a_2
X_5429_ VPWR VGND VPWR VGND _0862_ _0897_ _0876_ _0845_ _0898_ ZI_sky130_fd_sc_hd__or4_2
X_8148_ VGND VPWR _3523_ _2309_ _3043_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8079_ VGND VPWR VGND VPWR _0001_ _3751_ _4099_ _3461_ _3777_ ZI_sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_38_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_84_217 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_38_634 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_38_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_108_533 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_65_475 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_52_136 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_60_180 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4800_ VPWR VGND VGND VPWR _3906_ _0275_ _3974_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_28_133 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5780_ VPWR VGND VPWR VGND _0975_ _0841_ _0690_ _0710_ _1243_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_28_166 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_29_667 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4731_ VGND VPWR VGND VPWR _3978_ _3854_ _0207_ _4036_ ZI_sky130_fd_sc_hd__a21oi_2
X_4662_ VPWR VGND VPWR VGND _4174_ _4198_ _4186_ _4162_ _0139_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_83_272 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7450_ VPWR VGND _2888_ _2887_ _1677_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_56_486 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6401_ VPWR VGND VPWR VGND _1854_ _1858_ _1856_ _1853_ _1859_ ZI_sky130_fd_sc_hd__or4_2
X_7381_ VGND VPWR _2824_ _1061_ _2823_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_169 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_101_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4593_ VPWR VGND VPWR VGND _4129_ _4010_ _3926_ _3903_ _4005_ _4130_ ZI_sky130_fd_sc_hd__a221o_2
X_6332_ VGND VPWR VGND VPWR _1381_ _1344_ _1443_ _1791_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_101_73 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6263_ VPWR VGND VPWR VGND _1718_ _1722_ _1720_ _1715_ _1723_ ZI_sky130_fd_sc_hd__or4_2
X_8002_ VGND VPWR VPWR VGND _3389_ _3388_ _3391_ _3265_ _3390_ ZI_sky130_fd_sc_hd__o211a_2
X_5214_ VGND VPWR _0684_ _0586_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_86_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6194_ VPWR VGND VGND VPWR _1655_ _1389_ _1441_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_36_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5145_ VGND VPWR _0615_ _0614_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_98_309 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5076_ VGND VPWR _0546_ _0545_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5978_ VGND VPWR _1440_ _1409_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_19_100 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4929_ VPWR VGND VGND VPWR _0278_ _0176_ _3949_ _4019_ _3946_ _0402_ ZI_sky130_fd_sc_hd__a311o_2
X_7717_ VGND VPWR _3132_ _0377_ _0478_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_7648_ VPWR VGND VGND VPWR _3069_ _3066_ _3068_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_62_467 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7579_ VPWR VGND _3006_ block[115] round_key[115] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_15_372 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_62_489 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_106_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_57_228 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_31_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_38_464 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_25_103 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_26_648 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_25_147 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_80_253 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_80_275 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_21_331 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_80_297 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_0_225 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6950_ VGND VPWR VGND VPWR _2403_ _2302_ _2228_ _2119_ ZI_sky130_fd_sc_hd__o21a_2
X_5901_ VGND VPWR _1363_ _1362_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6881_ VGND VPWR VPWR VGND _2226_ _2333_ _2271_ _2334_ ZI_sky130_fd_sc_hd__or3_2
X_5832_ VGND VPWR VGND VPWR _0538_ _1290_ _1291_ _1292_ _1294_ _1293_ ZI_sky130_fd_sc_hd__o41ai_2
X_5763_ VGND VPWR VGND VPWR _1227_ _3756_ _1226_ _1204_ ZI_sky130_fd_sc_hd__o21a_2
X_7502_ VPWR VGND _2936_ block[12] round_key[12] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_84_581 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4714_ VPWR VGND VPWR VGND _0175_ _0189_ _0180_ _0172_ _0190_ ZI_sky130_fd_sc_hd__or4_2
X_8482_ VGND VPWR VPWR VGND clk _0084_ reset_n new_block[41] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_71_220 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5694_ VPWR VGND VPWR VGND _1159_ _0895_ _1158_ ZI_sky130_fd_sc_hd__or2_2
X_4645_ VGND VPWR VGND VPWR _4125_ _4181_ _3982_ _4178_ _4182_ ZI_sky130_fd_sc_hd__o22a_2
X_7433_ VGND VPWR VGND VPWR _2800_ new_block[70] _2872_ _2870_ _0475_ _0049_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_24_180 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7364_ VPWR VGND VPWR VGND _2797_ _2786_ _2808_ _2703_ _0241_ _2809_ ZI_sky130_fd_sc_hd__a221o_2
X_4576_ VPWR VGND VPWR VGND _3938_ _4112_ _4111_ _3922_ _4113_ ZI_sky130_fd_sc_hd__or4_2
X_6315_ VPWR VGND VPWR VGND _1308_ _1440_ _1491_ _1522_ _1774_ ZI_sky130_fd_sc_hd__a22o_2
X_7295_ VGND VPWR VPWR VGND _2741_ _2733_ _2743_ _1277_ _2742_ ZI_sky130_fd_sc_hd__o211a_2
X_6246_ VGND VPWR VGND VPWR _1704_ _1515_ _1705_ _1417_ _1706_ _1463_ ZI_sky130_fd_sc_hd__a2111o_2
X_6177_ VPWR VGND VPWR VGND _1635_ _1637_ _1636_ _1597_ _1638_ ZI_sky130_fd_sc_hd__or4_2
X_5128_ _0530_ _0598_ _3753_ _0576_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_99_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5059_ VPWR VGND VGND VPWR sword_ctr_reg\[0\] sword_ctr_reg\[1\] new_block[105] _0529_
+ ZI_sky130_fd_sc_hd__nor3_2
XFILLER_0_1_91 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_109_138 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_109_105 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_109_Right_109 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_23_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_62_253 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_30_161 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_26_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_301 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_45_209 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_389 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_1_501 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4430_ VGND VPWR VGND VPWR _3966_ _3965_ _3968_ _3967_ ZI_sky130_fd_sc_hd__a21oi_2
X_6100_ VGND VPWR VPWR VGND _1485_ _1561_ _1451_ _1562_ ZI_sky130_fd_sc_hd__or3_2
X_4361_ VGND VPWR VGND VPWR _3899_ _3898_ _3897_ _3893_ ZI_sky130_fd_sc_hd__o21a_2
X_7080_ VGND VPWR VGND VPWR _2531_ _2102_ _2256_ _2265_ ZI_sky130_fd_sc_hd__o21a_2
X_4292_ VPWR VGND VGND VPWR _3774_ _3827_ _3829_ _3830_ ZI_sky130_fd_sc_hd__nor3_2
XFILLER_0_67_44 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6031_ _1353_ _1493_ _1338_ _1363_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_7982_ VGND VPWR _3373_ _3371_ _3372_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_70 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_49_515 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6933_ _2060_ _2386_ _2099_ _2223_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_16_92 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6864_ VGND VPWR _2318_ _2315_ _2317_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_107_94 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5815_ VGND VPWR VPWR VGND _1275_ _1270_ _1278_ _1277_ _1276_ ZI_sky130_fd_sc_hd__o211a_2
X_6795_ VGND VPWR _2115_ _2168_ _2249_ _2236_ VPWR VGND ZI_sky130_fd_sc_hd__o21ai_2
XFILLER_0_107_609 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_17_445 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_44_220 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_8534_ VGND VPWR VPWR VGND clk _0136_ reset_n new_block[29] ZI_sky130_fd_sc_hd__dfrtp_2
X_5746_ VGND VPWR VGND VPWR _1209_ _0856_ _0652_ _1210_ ZI_sky130_fd_sc_hd__a21o_2
X_5677_ VGND VPWR VGND VPWR _1142_ _1130_ _1143_ _1001_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_44_253 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8465_ VGND VPWR VPWR VGND clk _0067_ reset_n new_block[88] ZI_sky130_fd_sc_hd__dfrtp_2
X_4628_ VGND VPWR VPWR VGND _3870_ _3998_ _3948_ _4165_ ZI_sky130_fd_sc_hd__or3_2
X_7416_ VGND VPWR _2857_ _4093_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_8396_ VPWR VGND VPWR VGND _3521_ _4093_ _3746_ _0169_ _1762_ _3747_ ZI_sky130_fd_sc_hd__a221o_2
X_7347_ VPWR VGND VGND VPWR _2793_ _2789_ _2792_ ZI_sky130_fd_sc_hd__nand2_2
X_4559_ VGND VPWR _4097_ _3822_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7278_ VPWR VGND VPWR VGND _2719_ _2725_ _2721_ _2654_ _2726_ ZI_sky130_fd_sc_hd__or4_2
X_6229_ VPWR VGND _1690_ _1689_ _1688_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_79_183 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_95_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_67_389 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_55_529 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_94_197 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_63_573 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5600_ VGND VPWR _1067_ _1063_ _1066_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6580_ VPWR VGND VPWR VGND _1788_ _1654_ _2035_ _2034_ _1716_ ZI_sky130_fd_sc_hd__or4b_2
XFILLER_0_6_637 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5531_ VGND VPWR _0999_ _0996_ _0998_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_253 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8250_ VPWR VGND _3615_ _2835_ _2790_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_112_601 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5462_ VPWR VGND VPWR VGND _0929_ _0841_ _0612_ _0711_ _0930_ ZI_sky130_fd_sc_hd__a22o_2
X_7201_ VPWR VGND VPWR VGND _2468_ _2222_ _2194_ _2073_ _2171_ _2650_ ZI_sky130_fd_sc_hd__a221o_2
X_4413_ _3945_ _3951_ _3949_ _3950_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8181_ VGND VPWR _3553_ _3551_ _3552_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_111_144 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_78_65 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5393_ VPWR VGND VPWR VGND _0849_ _0861_ _0858_ _0848_ _0862_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_1_386 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_10_632 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4344_ VPWR VGND VGND VPWR _3882_ _3878_ _3881_ ZI_sky130_fd_sc_hd__nand2_2
X_7132_ VGND VPWR VGND VPWR _2336_ _2299_ _2579_ _2580_ _2582_ _2581_ ZI_sky130_fd_sc_hd__a2111o_2
X_7063_ VGND VPWR VGND VPWR _2514_ _2196_ _2190_ _2512_ _2513_ ZI_sky130_fd_sc_hd__a211o_2
X_6014_ VPWR VGND VGND VPWR _1475_ _1476_ _1473_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_94_53 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4275_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[99] sword_ctr_reg\[0\] _3813_
+ ZI_sky130_fd_sc_hd__or3_2
X_7965_ VGND VPWR VGND VPWR _3331_ new_block[53] _3357_ _3354_ _1943_ _0096_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_49_301 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7896_ VGND VPWR VGND VPWR _3240_ new_block[47] _3294_ _3291_ _1268_ _0090_ ZI_sky130_fd_sc_hd__o32a_2
X_6916_ VPWR VGND VPWR VGND _2193_ _2368_ _2102_ _2235_ _2369_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_92_602 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_77_665 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6847_ VGND VPWR VGND VPWR _2301_ _2300_ _2168_ _2120_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_76_153 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6778_ VPWR VGND VPWR VGND _2155_ _2231_ _2229_ _2230_ _2232_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_92_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5729_ VGND VPWR _1194_ _0986_ _1193_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_573 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_8517_ VGND VPWR VPWR VGND clk _0119_ reset_n new_block[12] ZI_sky130_fd_sc_hd__dfrtp_2
X_8448_ VGND VPWR VPWR VGND clk _0050_ reset_n new_block[71] ZI_sky130_fd_sc_hd__dfrtp_2
X_8379_ VGND VPWR _3731_ _1563_ _1571_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_598 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_99_289 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_23_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_83_602 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_2_106 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_3_629 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_152 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_48_79 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_3_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Left_161 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4962_ VPWR VGND _0435_ _0153_ _4076_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7750_ VPWR VGND _3162_ _1760_ _1566_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6701_ VGND VPWR _2155_ _2154_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7681_ VGND VPWR _3099_ _0240_ _0309_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_473 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4893_ VPWR VGND _0367_ round_key[67] new_block[67] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6632_ sword_ctr_reg\[1\] _2086_ sword_ctr_reg\[0\] new_block[26] VPWR VGND VPWR
+ VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_27_573 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6563_ VPWR VGND VPWR VGND _1361_ _1464_ _1354_ _1376_ _2018_ ZI_sky130_fd_sc_hd__a22o_2
X_8302_ VGND VPWR _3662_ _0808_ _1068_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5514_ VPWR VGND VPWR VGND _0974_ _0981_ _0977_ _0972_ _0982_ ZI_sky130_fd_sc_hd__or4_2
X_6494_ VPWR VGND _1951_ _1898_ _1578_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_57_Left_170 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_14_289 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5445_ VGND VPWR _0914_ _0911_ _0913_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8233_ VPWR VGND VGND VPWR _3600_ _3596_ _3599_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_1_150 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8164_ VGND VPWR VPWR VGND _3536_ _3535_ _3538_ _3448_ _3537_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_66_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7115_ VPWR VGND VPWR VGND _4100_ _1909_ _2565_ _1959_ _2564_ _2566_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_100_637 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5376_ VPWR VGND VGND VPWR _0836_ _0840_ _0844_ _0845_ ZI_sky130_fd_sc_hd__nor3_2
X_8095_ VGND VPWR _3475_ _4087_ _1586_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4327_ VGND VPWR _3865_ _3864_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_4258_ VGND VPWR _3796_ _3787_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7046_ VPWR VGND VPWR VGND _4100_ _1909_ _2497_ _1959_ _2496_ _2498_ ZI_sky130_fd_sc_hd__a221o_2
X_7948_ VPWR VGND _3342_ block[84] round_key[84] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_49_120 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_9_261 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7879_ VGND VPWR _3279_ _2547_ _3278_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_134 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_80_638 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_16_Right_16 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_68_473 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_95_270 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_55_178 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_25_Right_25 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_70_159 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_70_148 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_51_362 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5230_ VPWR VGND _0608_ _0700_ _0586_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5161_ VGND VPWR VPWR VGND _0537_ _0543_ _3774_ _0631_ ZI_sky130_fd_sc_hd__or3_2
X_5092_ VGND VPWR VGND VPWR _0538_ _0558_ _0559_ _0560_ _0562_ _0561_ ZI_sky130_fd_sc_hd__o41ai_2
XPHY_EDGE_ROW_34_Right_34 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5994_ VPWR VGND VGND VPWR _1436_ _1456_ _1455_ ZI_sky130_fd_sc_hd__nor2_2
X_7802_ VPWR VGND VPWR VGND _3150_ _3159_ _3209_ _3139_ _0907_ _3210_ ZI_sky130_fd_sc_hd__a221o_2
X_4945_ VPWR VGND VPWR VGND _4042_ _4031_ _3997_ _0185_ _0418_ ZI_sky130_fd_sc_hd__a22o_2
X_7733_ VGND VPWR VGND VPWR _3147_ _3146_ _3145_ _3143_ ZI_sky130_fd_sc_hd__o21a_2
X_7664_ VGND VPWR _3083_ _0145_ _0310_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4876_ VPWR VGND VPWR VGND _3950_ _3926_ _3911_ _4012_ _0350_ ZI_sky130_fd_sc_hd__a22o_2
X_7595_ VPWR VGND _3020_ _2497_ _2313_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_43_Right_43 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_46_178 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6615_ VGND VPWR VGND VPWR _0538_ _2065_ _2066_ _2067_ _2069_ _2068_ ZI_sky130_fd_sc_hd__o41ai_2
X_6546_ VGND VPWR _2002_ _2000_ _2001_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_587 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_70_660 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6477_ VGND VPWR VGND VPWR _1385_ _1357_ _1934_ _1653_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_30_557 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5428_ VPWR VGND VPWR VGND _0882_ _0896_ _0890_ _0733_ _0897_ ZI_sky130_fd_sc_hd__or4_2
X_8216_ VPWR VGND VPWR VGND _3575_ _3490_ _3584_ _3583_ _1578_ _3585_ ZI_sky130_fd_sc_hd__a221o_2
X_8147_ VGND VPWR VGND VPWR _3462_ new_block[6] _3522_ _3517_ _0475_ _0113_ ZI_sky130_fd_sc_hd__o32a_2
X_5359_ VGND VPWR VGND VPWR _0828_ _0684_ _0592_ _0609_ _0532_ ZI_sky130_fd_sc_hd__and4_2
X_8078_ VPWR VGND VPWR VGND _3459_ _3367_ _3457_ _3328_ _1566_ _3460_ ZI_sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_52_Right_52 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7029_ VPWR VGND VGND VPWR _2480_ _2479_ _2073_ _2219_ _2229_ _2481_ ZI_sky130_fd_sc_hd__a311o_2
XFILLER_0_97_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_38_613 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_84_229 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_38_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_65_410 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_53_605 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_61_Right_61 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_108_545 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_108_589 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_110_209 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_60_192 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_29_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_45_69 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_61_24 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_61_57 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4730_ VGND VPWR VGND VPWR _4168_ _3845_ _3988_ _3874_ _0206_ ZI_sky130_fd_sc_hd__a2bb2o_2
X_4661_ VPWR VGND VPWR VGND _4194_ _4034_ _4196_ _4197_ _4198_ ZI_sky130_fd_sc_hd__or4bb_2
XFILLER_0_56_498 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7380_ VPWR VGND _2823_ _1138_ _1135_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6400_ VGND VPWR VGND VPWR _1857_ _1319_ _1346_ _1414_ _1858_ ZI_sky130_fd_sc_hd__a31o_2
X_6331_ VGND VPWR VPWR VGND _1787_ _1789_ _1784_ _1790_ ZI_sky130_fd_sc_hd__or3_2
X_4592_ VPWR VGND VGND VPWR _3887_ _4129_ _3854_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_10_61 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_101_85 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6262_ VPWR VGND VPWR VGND _1721_ _1389_ _1432_ _1308_ _1332_ _1722_ ZI_sky130_fd_sc_hd__a221o_2
X_8001_ VPWR VGND VGND VPWR _3390_ _3388_ _3389_ ZI_sky130_fd_sc_hd__nand2_2
X_6193_ VGND VPWR VGND VPWR _1535_ _1371_ _1653_ _1654_ ZI_sky130_fd_sc_hd__a21o_2
X_5213_ VPWR VGND VGND VPWR _0650_ _0683_ _0617_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_86_65 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5144_ VPWR VGND _0605_ _0614_ _0608_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_19_81 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5075_ VGND VPWR _0545_ _0544_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_29_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_79_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5977_ VPWR VGND VPWR VGND _1438_ _1434_ _1431_ _1432_ _1439_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_47_421 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7716_ VGND VPWR VGND VPWR _2799_ new_block[94] _3131_ _3129_ _2731_ _0073_ ZI_sky130_fd_sc_hd__o32a_2
X_4928_ VGND VPWR VGND VPWR _0400_ _3948_ _3945_ _4134_ _0401_ ZI_sky130_fd_sc_hd__a31o_2
XFILLER_0_34_115 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_47_487 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7647_ VGND VPWR _3068_ _0370_ _3067_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4859_ VGND VPWR VGND VPWR _0333_ _0332_ _0330_ _0328_ _0326_ ZI_sky130_fd_sc_hd__and4_2
X_7578_ VGND VPWR VPWR VGND _3003_ _2998_ _3005_ _2855_ _3004_ ZI_sky130_fd_sc_hd__o211a_2
X_6529_ VPWR VGND _1349_ _1985_ _1512_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
XFILLER_0_100_220 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_100_253 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_100_264 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_15_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_549 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_31_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_80_243 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_80_232 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_80_265 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_0_237 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_104_581 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5900_ VGND VPWR VPWR VGND _1316_ _1317_ _3832_ _1362_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_88_332 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6880_ VPWR VGND VPWR VGND _2186_ _2300_ _2135_ _2265_ _2333_ ZI_sky130_fd_sc_hd__a22o_2
X_5831_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[113] sword_ctr_reg\[0\] _1293_
+ ZI_sky130_fd_sc_hd__or3_2
X_5762_ VPWR VGND VPWR VGND _0845_ _1225_ _1213_ _0720_ _1226_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_16_104 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7501_ VGND VPWR VPWR VGND _2933_ _2931_ _2935_ _2855_ _2934_ ZI_sky130_fd_sc_hd__o211a_2
X_4713_ VPWR VGND VPWR VGND _0188_ _0189_ _0184_ _0187_ ZI_sky130_fd_sc_hd__or3b_2
X_8481_ VGND VPWR VPWR VGND clk _0083_ reset_n new_block[40] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_137 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_44_435 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5693_ VPWR VGND VPWR VGND _0833_ _0613_ _0712_ _0662_ _0710_ _1158_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_21_71 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4644_ VGND VPWR _4181_ _3992_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7432_ VPWR VGND VPWR VGND _2797_ _2871_ _2857_ _2703_ _4067_ _2872_ ZI_sky130_fd_sc_hd__a221o_2
X_4575_ VGND VPWR VGND VPWR _3903_ _3900_ _4047_ _4112_ ZI_sky130_fd_sc_hd__a21o_2
X_7363_ VPWR VGND _2808_ block[33] round_key[33] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6314_ VGND VPWR VGND VPWR _1332_ _1491_ _1550_ _1773_ ZI_sky130_fd_sc_hd__a21o_2
XFILLER_0_40_641 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7294_ VPWR VGND VGND VPWR _2742_ _2733_ _2741_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_12_365 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6245_ VGND VPWR VGND VPWR _1535_ _1371_ _1705_ _1384_ ZI_sky130_fd_sc_hd__a21oi_2
X_6176_ VPWR VGND VGND VPWR _1416_ _1637_ _1370_ ZI_sky130_fd_sc_hd__nor2_2
X_5127_ VPWR VGND VPWR VGND _0545_ _0596_ _0592_ _0595_ _0597_ ZI_sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_2_Right_2 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5058_ VGND VPWR VGND VPWR sword_ctr_reg\[1\] sword_ctr_reg\[0\] new_block[73] _0528_
+ ZI_sky130_fd_sc_hd__nand3b_2
XFILLER_0_98_107 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_94_346 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_105_389 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_101_551 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Left_124 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_66_560 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_26_468 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_41_416 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_81_574 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_20_Left_133 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_41_427 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_41_449 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_6_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4360_ VGND VPWR _3898_ _3878_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_1_557 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_111_337 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4291_ VPWR VGND VGND VPWR _3828_ _3829_ new_block[101] ZI_sky130_fd_sc_hd__nor2_2
X_6030_ VPWR VGND VPWR VGND _1491_ _1489_ _1426_ _1428_ _1492_ ZI_sky130_fd_sc_hd__a22o_2
X_7981_ VPWR VGND _3372_ _4074_ _4068_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_107_51 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_89_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6932_ VGND VPWR VGND VPWR _2385_ _2147_ _2297_ _2207_ _2327_ ZI_sky130_fd_sc_hd__and4_2
X_6863_ VGND VPWR _2317_ _2048_ _2316_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5814_ VGND VPWR _1277_ _0365_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_8_123 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6794_ VPWR VGND VGND VPWR _2144_ _2248_ _2097_ ZI_sky130_fd_sc_hd__nor2_2
X_8533_ VGND VPWR VPWR VGND clk _0135_ reset_n new_block[28] ZI_sky130_fd_sc_hd__dfrtp_2
X_5745_ VPWR VGND VGND VPWR _1209_ _0684_ _0626_ ZI_sky130_fd_sc_hd__nand2_2
X_5676_ VGND VPWR _1142_ _1134_ _1141_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8464_ VGND VPWR VPWR VGND clk _0066_ reset_n new_block[87] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_340 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7415_ VGND VPWR VPWR VGND _2853_ _2847_ _2856_ _2855_ _2854_ ZI_sky130_fd_sc_hd__o211a_2
XFILLER_0_32_449 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_44_287 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_4627_ VPWR VGND VPWR VGND _4164_ _3971_ _3988_ ZI_sky130_fd_sc_hd__or2_2
XFILLER_0_13_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8395_ VPWR VGND _3746_ block[31] round_key[31] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_7346_ VGND VPWR _2792_ _2790_ _2791_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4558_ VPWR VGND VPWR VGND _4096_ round_key[64] block[64] ZI_sky130_fd_sc_hd__or2_2
X_4489_ VPWR VGND VGND VPWR _4026_ _4024_ _4008_ _3913_ _4019_ _4027_ ZI_sky130_fd_sc_hd__a311o_2
X_7277_ VPWR VGND VPWR VGND _2722_ _2724_ _2723_ _2433_ _2725_ ZI_sky130_fd_sc_hd__or4_2
X_6228_ VPWR VGND _1689_ round_key[14] new_block[14] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6159_ VGND VPWR VGND VPWR _1620_ _1341_ _1523_ _1619_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_82_305 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_63_585 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_31_471 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_101_370 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_5_126 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5530_ VPWR VGND _0998_ _0997_ _0800_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_26_265 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5461_ VPWR VGND _0630_ _0929_ _0705_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_7200_ VGND VPWR VGND VPWR _2649_ _2219_ _2648_ _2381_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_112_613 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_4412_ _3891_ _3950_ _3831_ _3892_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
X_8180_ VGND VPWR _3552_ _0306_ _3076_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_657 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5392_ VPWR VGND VPWR VGND _0860_ _0787_ _0859_ _0675_ _0702_ _0861_ ZI_sky130_fd_sc_hd__a221o_2
X_4343_ VPWR VGND VGND VPWR _3880_ _3881_ _3809_ _3814_ ZI_sky130_fd_sc_hd__nor3b_2
XPHY_EDGE_ROW_99_Right_99 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_7131_ VPWR VGND VPWR VGND _2265_ _2158_ _2327_ _2216_ _2581_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_78_77 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7062_ VPWR VGND VPWR VGND _2345_ _2279_ _2260_ _2154_ _2513_ ZI_sky130_fd_sc_hd__a22o_2
X_4274_ VGND VPWR VPWR VGND sword_ctr_reg\[0\] _3812_ new_block[35] ZI_sky130_fd_sc_hd__and2b_2
X_6013_ VPWR VGND VGND VPWR _1475_ _1474_ _1375_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_94_65 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7964_ VGND VPWR VGND VPWR _3357_ _3355_ _4094_ _3356_ _3150_ ZI_sky130_fd_sc_hd__a211o_2
XFILLER_0_11_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_49_324 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6915_ VGND VPWR _2368_ _2281_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7895_ VPWR VGND VPWR VGND _3219_ _3257_ _3293_ _3237_ _3292_ _3294_ ZI_sky130_fd_sc_hd__a221o_2
XFILLER_0_92_614 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6846_ VGND VPWR _2300_ _2267_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_76_176 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_76_165 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6777_ VGND VPWR _2231_ _2204_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5728_ VGND VPWR _1193_ _1132_ _1192_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8516_ VGND VPWR VPWR VGND clk _0118_ reset_n new_block[11] ZI_sky130_fd_sc_hd__dfrtp_2
X_8447_ VGND VPWR VPWR VGND clk _0049_ reset_n new_block[70] ZI_sky130_fd_sc_hd__dfrtp_2
X_5659_ VGND VPWR VGND VPWR _1125_ _3756_ _1124_ _1098_ ZI_sky130_fd_sc_hd__o21a_2
X_8378_ VGND VPWR VGND VPWR _3640_ new_block[29] _3730_ _3728_ _2686_ _0136_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_40_290 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7329_ VPWR VGND _2776_ _2309_ _2011_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_7_91 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_99_202 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_99_246 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_99_268 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_67_121 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_23_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_67_176 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_67_165 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_82_157 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_23_257 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_64_57 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_98_290 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4961_ VGND VPWR _0434_ _0230_ _0231_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4892_ VGND VPWR _0366_ _0365_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7680_ VGND VPWR _3098_ _0301_ _0375_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6700_ VPWR VGND VGND VPWR _2147_ _2154_ _2095_ ZI_sky130_fd_sc_hd__nor2_2
X_6631_ VGND VPWR VGND VPWR _2085_ sword_ctr_reg\[0\] new_block[90] sword_ctr_reg\[1\]
+ ZI_sky130_fd_sc_hd__and3b_2
XFILLER_0_104_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_13_83 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_104_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8301_ VGND VPWR _3661_ _1273_ _3660_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6562_ VGND VPWR VPWR VGND _2017_ _1346_ _1351_ _1464_ _1341_ ZI_sky130_fd_sc_hd__o31a_2
XFILLER_0_14_235 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_5513_ VPWR VGND VPWR VGND _0790_ _0980_ _0979_ _0978_ _0981_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_42_533 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6493_ VGND VPWR _1950_ _1680_ _1949_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_5444_ VGND VPWR _0913_ _0808_ _0912_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_577 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_8232_ VGND VPWR _3599_ _3597_ _3598_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_8163_ VPWR VGND VGND VPWR _3537_ _3535_ _3536_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_1_162 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_7114_ VPWR VGND _2565_ new_block[123] round_key[123] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5375_ VPWR VGND VPWR VGND _0844_ _0842_ _0843_ ZI_sky130_fd_sc_hd__or2_2
XFILLER_0_59_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_1_195 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8094_ VGND VPWR _3474_ _1770_ _2311_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_4326_ VPWR VGND VPWR VGND _3863_ _3847_ _3824_ _3830_ _3864_ ZI_sky130_fd_sc_hd__or4_2
X_7045_ VPWR VGND _2497_ new_block[122] round_key[122] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_4257_ VGND VPWR _3795_ _3794_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7947_ VGND VPWR VGND VPWR _3341_ _3340_ _3338_ _3332_ ZI_sky130_fd_sc_hd__o21a_2
X_7878_ VGND VPWR _3278_ _1198_ _2011_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_143 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_6829_ VGND VPWR VGND VPWR _2283_ _2282_ _2279_ _2190_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_18_596 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_33_544 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_13_290 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_0_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_34_16 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_71_617 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_24_522 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_51_374 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_106_281 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_59_57 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5160_ VGND VPWR _0630_ _0629_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5091_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[110] sword_ctr_reg\[0\] _0561_
+ ZI_sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_3_Left_116 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5993_ VGND VPWR VGND VPWR _1294_ _1347_ _1455_ _3796_ ZI_sky130_fd_sc_hd__a21oi_2
X_7801_ VPWR VGND _3209_ block[6] round_key[6] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_59_441 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_91_88 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7732_ VGND VPWR VGND VPWR _3145_ _3143_ _3146_ _3028_ ZI_sky130_fd_sc_hd__a21oi_2
X_4944_ VPWR VGND VPWR VGND _0403_ _0416_ _0411_ _0398_ _0417_ ZI_sky130_fd_sc_hd__or4_2
X_7663_ VGND VPWR VGND VPWR new_block[90] _2800_ _2483_ _3082_ _0069_ ZI_sky130_fd_sc_hd__o22a_2
X_4875_ VPWR VGND VPWR VGND _0349_ _0343_ _0348_ ZI_sky130_fd_sc_hd__or2_2
XFILLER_0_62_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7594_ VGND VPWR VGND VPWR new_block[84] _2800_ _1884_ _3019_ _0063_ ZI_sky130_fd_sc_hd__o22a_2
X_6614_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] new_block[127] sword_ctr_reg\[0\] _2068_
+ ZI_sky130_fd_sc_hd__or3_2
X_6545_ VGND VPWR _2001_ _1569_ _1680_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_599 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_6476_ VGND VPWR VGND VPWR _1932_ _1395_ _1521_ _1529_ _1933_ ZI_sky130_fd_sc_hd__a31o_2
X_8215_ VPWR VGND _3584_ block[77] round_key[77] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_30_569 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5427_ VPWR VGND VPWR VGND _0893_ _0895_ _0894_ _0892_ _0896_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_100_402 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5358_ VPWR VGND VGND VPWR _0827_ _3755_ _0590_ ZI_sky130_fd_sc_hd__nand2_2
X_8146_ VPWR VGND VGND VPWR _3521_ _3520_ _0162_ _3518_ _3519_ _3522_ ZI_sky130_fd_sc_hd__a311o_2
X_4309_ VPWR VGND _3753_ _3847_ _3843_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_8077_ VGND VPWR _3459_ _3458_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5289_ VGND VPWR VGND VPWR _0756_ _0748_ _0758_ _0759_ ZI_sky130_fd_sc_hd__a21o_2
X_7028_ _2339_ _2480_ _2187_ _2246_ VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__and3_2
XFILLER_0_37_102 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_37_124 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_65_422 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_108_502 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_108_557 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_33_374 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_29_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_189 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_85_Left_198 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_56_466 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_9_15 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4660_ VGND VPWR VGND VPWR _3895_ _3896_ _4116_ _3906_ _4197_ ZI_sky130_fd_sc_hd__o22a_2
XFILLER_0_56_477 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_83_296 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_6330_ VGND VPWR VGND VPWR _1789_ _1529_ _1337_ _1741_ _1788_ ZI_sky130_fd_sc_hd__a211o_2
X_4591_ VPWR VGND VPWR VGND _4127_ _4128_ _4124_ _4126_ ZI_sky130_fd_sc_hd__or3b_2
X_6261_ VPWR VGND _1613_ _1721_ _1639_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_8000_ VGND VPWR _3389_ _0914_ _1131_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6192_ VGND VPWR _1653_ _1652_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5212_ VPWR VGND _0634_ _0682_ _0670_ VPWR VGND ZI_sky130_fd_sc_hd__and2_2
X_5143_ VGND VPWR _0613_ _0612_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_86_77 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5074_ VPWR VGND VGND VPWR _3796_ _0537_ _0543_ _0544_ ZI_sky130_fd_sc_hd__nor3_2
XFILLER_0_35_81 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_5976_ VGND VPWR _1438_ _1437_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_47_444 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7715_ VPWR VGND VPWR VGND _2995_ _2960_ _3130_ _2984_ _0142_ _3131_ ZI_sky130_fd_sc_hd__a221o_2
X_4927_ VGND VPWR VGND VPWR _4052_ _3882_ _0400_ _3987_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_34_105 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4858_ VPWR VGND VGND VPWR _4153_ _3896_ _4175_ _3906_ _0332_ _0331_ ZI_sky130_fd_sc_hd__o221a_2
X_7646_ VGND VPWR _3067_ _4064_ _0298_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_127 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_105_505 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7577_ VPWR VGND VGND VPWR _3004_ _2998_ _3003_ ZI_sky130_fd_sc_hd__nand2_2
X_4789_ VPWR VGND VPWR VGND _0259_ _0263_ _0260_ _4137_ _0264_ ZI_sky130_fd_sc_hd__or4_2
X_6528_ VGND VPWR VGND VPWR _1984_ _1534_ _1632_ _1727_ ZI_sky130_fd_sc_hd__o21a_2
X_6459_ VPWR VGND VPWR VGND _1913_ _1915_ _1914_ _1912_ _1916_ ZI_sky130_fd_sc_hd__or4_2
X_8129_ VGND VPWR VGND VPWR _3505_ _3504_ _3506_ _3339_ ZI_sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_388 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_38_433 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_31_39 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_93_583 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_108_365 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_40_108 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_33_160 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_0_249 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_93_Left_206 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5830_ VGND VPWR VPWR VGND sword_ctr_reg\[1\] _1292_ new_block[81] ZI_sky130_fd_sc_hd__and2b_2
XFILLER_0_69_591 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_8_305 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5761_ VPWR VGND VPWR VGND _1031_ _1224_ _1217_ _0821_ _1225_ ZI_sky130_fd_sc_hd__or4_2
XFILLER_0_17_606 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_17_617 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7500_ VPWR VGND VGND VPWR _2934_ _2931_ _2933_ ZI_sky130_fd_sc_hd__nand2_2
X_8480_ VGND VPWR VPWR VGND clk _0082_ reset_n new_block[39] ZI_sky130_fd_sc_hd__dfrtp_2
X_4712_ VGND VPWR VGND VPWR _3935_ _3949_ _3998_ _3930_ _3967_ _0188_ ZI_sky130_fd_sc_hd__o32a_2
XFILLER_0_44_447 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_112_41 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7431_ VPWR VGND _2871_ block[38] round_key[38] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5692_ VGND VPWR VGND VPWR _1157_ _0722_ _0776_ _0646_ ZI_sky130_fd_sc_hd__o21a_2
XFILLER_0_4_522 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_4643_ VPWR VGND VGND VPWR _4052_ _3906_ _4131_ _3921_ _4180_ _4179_ ZI_sky130_fd_sc_hd__o221a_2
XFILLER_0_112_85 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_21_83 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
X_7362_ VGND VPWR VPWR VGND _2805_ _0797_ _2807_ _1277_ _2806_ ZI_sky130_fd_sc_hd__o211a_2
X_4574_ VPWR VGND VGND VPWR _4110_ _4111_ _3984_ ZI_sky130_fd_sc_hd__nor2_2
X_6313_ VPWR VGND VPWR VGND _1521_ _1395_ _1434_ _1522_ _1619_ _1772_ ZI_sky130_fd_sc_hd__a221o_2
X_7293_ VGND VPWR _2741_ _2737_ _2740_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
X_6244_ VPWR VGND VGND VPWR _1653_ _1704_ _1357_ ZI_sky130_fd_sc_hd__nor2_2
X_6175_ VPWR VGND VGND VPWR _1405_ _1636_ _1307_ ZI_sky130_fd_sc_hd__nor2_2
X_5126_ VGND VPWR VGND VPWR _0576_ _0593_ _3880_ _0596_ ZI_sky130_fd_sc_hd__a21o_2
X_5057_ VGND VPWR VGND VPWR sword_ctr_reg\[0\] new_block[41] sword_ctr_reg\[1\] _0527_
+ ZI_sky130_fd_sc_hd__nand3b_2
XFILLER_0_79_333 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_5959_ VGND VPWR _1421_ _1420_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_90_520 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
XFILLER_0_7_393 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_7629_ VPWR VGND VGND VPWR _0149_ _3052_ _4090_ ZI_sky130_fd_sc_hd__nor2_2
XFILLER_0_30_141 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_101_574 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_98_631 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_85_325 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_38_274 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_109_641 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_66_572 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4290_ VGND VPWR _3828_ _3822_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7980_ VPWR VGND _3371_ _3133_ _0373_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
XFILLER_0_89_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_88_141 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6931_ VPWR VGND VPWR VGND _2380_ _2383_ _2381_ _2379_ _2384_ ZI_sky130_fd_sc_hd__or4_2
X_6862_ VPWR VGND _2316_ _1961_ _1586_ VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_5813_ VPWR VGND VGND VPWR _1276_ _1270_ _1275_ ZI_sky130_fd_sc_hd__nand2_2
XFILLER_0_8_135 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_6793_ VPWR VGND VPWR VGND _2155_ _2246_ _2097_ _2233_ _2247_ ZI_sky130_fd_sc_hd__a22o_2
X_8532_ VGND VPWR VPWR VGND clk _0134_ reset_n new_block[27] ZI_sky130_fd_sc_hd__dfrtp_2
XFILLER_0_84_391 VGND VPWR VPWR VGND ZI_sky130_fd_sc_hd__decap_4
X_5744_ VPWR VGND VGND VPWR _1208_ _0628_ _0729_ ZI_sky130_fd_sc_hd__nand2_2
X_5675_ VGND VPWR _1141_ _1136_ _1140_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_458 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
X_8463_ VGND VPWR VPWR VGND clk _0065_ reset_n new_block[86] ZI_sky130_fd_sc_hd__dfrtp_2
X_7414_ VGND VPWR _2855_ _0365_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
XFILLER_0_89_3 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_8394_ VGND VPWR VPWR VGND _3743_ _3742_ _3745_ _0366_ _3744_ ZI_sky130_fd_sc_hd__o211a_2
X_4626_ VPWR VGND VPWR VGND _3824_ _3895_ _3847_ _3890_ _4163_ ZI_sky130_fd_sc_hd__or4_2
X_7345_ VGND VPWR _2791_ _0912_ _1192_ VPWR VGND ZI_sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_653 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_4557_ VPWR VGND VGND VPWR _4095_ round_key[64] block[64] ZI_sky130_fd_sc_hd__nand2_2
X_4488_ VGND VPWR VGND VPWR _4025_ _3954_ _4026_ _3999_ ZI_sky130_fd_sc_hd__a21oi_2
X_7276_ VPWR VGND VPWR VGND _2237_ _2114_ _2216_ _2102_ _2131_ _2724_ ZI_sky130_fd_sc_hd__a221o_2
X_6227_ VPWR VGND _1688_ round_key[9] new_block[9] VPWR VGND ZI_sky130_fd_sc_hd__xor2_2
X_6158_ VPWR VGND VGND VPWR _1436_ _1619_ _1295_ ZI_sky130_fd_sc_hd__nor2_2
X_5109_ VGND VPWR _0579_ _0578_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_6089_ VGND VPWR VPWR VGND _1313_ _1318_ _1382_ _1551_ ZI_sky130_fd_sc_hd__or3_2
XFILLER_0_63_597 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_31_483 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_3
XFILLER_0_37_27 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_101_393 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
XFILLER_0_86_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
XFILLER_0_39_561 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_6
X_5460_ VGND VPWR VGND VPWR _0927_ _0923_ _0928_ _0924_ ZI_sky130_fd_sc_hd__a21bo_2
XFILLER_0_54_597 VPWR VGND VPWR VGND ZI_sky130_fd_sc_hd__decap_8
XFILLER_0_41_225 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_4411_ VGND VPWR _3949_ _3948_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_5391_ VPWR VGND VPWR VGND _0740_ _0741_ _0675_ _0669_ _0860_ ZI_sky130_fd_sc_hd__a22o_2
XFILLER_0_10_645 VGND VPWR VPWR VGND ZI_sky130_ef_sc_hd__decap_12
X_7130_ VGND VPWR VGND VPWR _2580_ _2208_ _2193_ _2112_ ZI_sky130_fd_sc_hd__o21a_2
X_4342_ VGND VPWR _3880_ _3879_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
X_7061_ VPWR VGND VPWR VGND _2144_ _2373_ _2112_ _2231_ _2512_ ZI_sky130_fd_sc_hd__a22o_2
X_4273_ sword_ctr_reg\[1\] _3811_ sword_ctr_reg\[0\] new_block[3] VPWR VGND VPWR VGND
+ ZI_sky130_fd_sc_hd__and3_2
X_6012_ VGND VPWR _1474_ _1369_ VPWR VGND ZI_sky130_fd_sc_hd__buf_1
.ends

.subckt sky130_fd_sc_hd__nor3_2 VPB VNB VGND VPWR A B C Y
X0 Y C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X6 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X10 a_281_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4bb_2 VNB VPB VGND VPWR A_N X C D B_N
X0 a_174_21# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1 a_174_21# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.33075 ps=1.705 w=0.42 l=0.15
X2 a_476_47# a_27_47# a_174_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33075 pd=1.705 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X5 a_548_47# a_505_280# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8 VPWR D a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND D a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 VPWR a_505_280# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X11 a_505_280# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X12 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_505_280# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X14 a_639_47# C a_548_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X15 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4_2 VNB VPB VGND VPWR B D Y A C
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_475_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y D a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12 a_475_297# C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_281_297# C a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X14 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X15 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_2 VNB VPB VGND VPWR X D C B A
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.27995 ps=1.615 w=1 l=0.15
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.06195 ps=0.715 w=0.42 l=0.15
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.17515 ps=1.265 w=0.65 l=0.15
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.07455 ps=0.775 w=0.42 l=0.15
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_2 VNB VPB VGND VPWR B1 B2 A2_N A1_N X
X0 VPWR a_82_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.435 as=0.135 ps=1.27 w=1 l=0.15
X1 a_646_47# B2 a_82_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_574_369# a_313_47# a_82_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0976 pd=0.945 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 a_574_369# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4 VGND a_82_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR B2 a_574_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0976 ps=0.945 w=0.64 l=0.15
X6 X a_82_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 X a_82_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8 a_313_47# A2_N a_313_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.0672 ps=0.85 w=0.64 l=0.15
X9 a_313_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X10 a_313_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.186 ps=1.435 w=0.64 l=0.15
X11 VGND A2_N a_313_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14175 pd=1.095 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_82_21# a_313_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.14175 ps=1.095 w=0.42 l=0.15
X13 VGND B1 a_646_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_2 VNB VPB VGND VPWR Y B1 A2 A1 C1
X0 a_286_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2 a_286_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X3 Y A2 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 VGND A1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X6 VGND A2 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 a_487_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_27_47# B1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR A1 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X13 a_487_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14 a_286_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22ai_2 VPB VNB VGND VPWR A1 A2 Y B2 B1
X0 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_475_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR A1 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.26975 pd=1.48 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12 a_475_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 Y A2 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X14 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.26975 ps=1.48 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_2 VNB VPB VGND VPWR B1 B2 A3 A2 A1 X
X0 a_429_297# A2 a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND A2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_345_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13975 ps=1.08 w=0.65 l=0.15
X5 a_345_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=1.61 w=1 l=0.15
X6 a_629_297# B2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR B1 a_629_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.19 ps=1.38 w=1 l=0.15
X8 a_79_21# B2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_345_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.1235 ps=1.03 w=0.65 l=0.15
X10 a_79_21# A3 a_429_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_345_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.26 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_2 VNB VPB VGND VPWR B1_N Y A2 A1
X0 a_397_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR B1_N a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 Y A2 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VGND A2 a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VGND A1 a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_28_297# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 Y a_28_297# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR a_28_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_397_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X9 a_229_47# a_28_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y a_28_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X11 a_229_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_229_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VPWR A1 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfstp_2 VPB VNB VPWR VGND Q SET_B D CLK
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.06705 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_1136_413# a_193_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X3 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06705 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X5 a_1228_47# a_27_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X6 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X8 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12495 pd=1.175 as=0.2184 ps=2.2 w=0.84 l=0.15
X10 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X11 VPWR a_1602_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1028_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VGND a_1602_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_1028_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.12495 ps=1.175 w=0.42 l=0.15
X18 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1028_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X20 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X21 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_1028_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0441 ps=0.63 w=0.42 l=0.15
X23 VPWR a_1178_261# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X24 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 a_1178_261# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2226 pd=2.21 as=0.12075 ps=1.165 w=0.84 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_1300_47# a_1178_261# a_1228_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X28 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X29 a_1178_261# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1404 pd=1.6 as=0.1137 ps=1.01 w=0.54 l=0.15
X30 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X31 VPWR SET_B a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12075 pd=1.165 as=0.1092 ps=1.36 w=0.42 l=0.15
X32 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X33 VGND SET_B a_1300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1137 pd=1.01 as=0.0441 ps=0.63 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32oi_2 VNB VPB VGND VPWR B2 B1 Y A1 A2 A3
X0 Y A1 a_478_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.3775 ps=1.755 w=1 l=0.15
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.305 ps=1.61 w=1 l=0.15
X3 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.335 ps=1.67 w=1 l=0.15
X4 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.1375 ps=1.275 w=1 l=0.15
X5 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3775 pd=1.755 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_478_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_478_47# A2 a_730_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND A3 a_730_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12025 ps=1.02 w=0.65 l=0.15
X10 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_730_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.20475 ps=1.93 w=0.65 l=0.15
X16 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.15 ps=1.3 w=1 l=0.15
X18 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X19 a_730_47# A2 a_478_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111oi_2 VNB VPB VGND VPWR A1 A2 D1 C1 B1 Y
X0 a_467_297# B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X1 a_287_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR A2 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X3 a_923_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.112125 ps=0.995 w=0.65 l=0.15
X4 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X5 a_28_297# B1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X7 a_28_297# C1 a_287_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X8 Y A1 a_923_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND A2 a_684_47# VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17875 ps=1.2 w=0.65 l=0.15
X10 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.105625 ps=0.975 w=0.65 l=0.15
X12 Y D1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_467_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=2.67 as=0.16 ps=1.32 w=1 l=0.15
X14 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.12675 ps=1.04 w=0.65 l=0.15
X16 VPWR A1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X17 a_115_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X18 a_467_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 a_684_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.2 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32o_2 VNB VPB VGND VPWR X A3 A2 B2 B1 A1
X0 VPWR A3 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X2 a_352_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.209625 ps=1.295 w=0.65 l=0.15
X3 a_549_47# A1 a_21_199# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 X a_21_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_21_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.209625 pd=1.295 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13975 ps=1.08 w=0.65 l=0.15
X7 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X8 a_299_297# B1 a_21_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_21_199# B2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND A3 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR a_21_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 X a_21_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_21_199# B1 a_352_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.115375 ps=1.005 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221ai_2 VNB VPB VGND VPWR Y B1 B2 A2 A1 C1
X0 Y A2 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_300_47# B2 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 a_300_47# B1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_300_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_734_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X7 a_28_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y C1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR B1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X11 a_382_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_28_47# B1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_28_47# B2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X15 Y B2 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VPWR A1 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND A2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_382_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X19 a_734_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_2 VPWR VGND VPB VNB B2 B1 Y A1 A2
X0 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_467_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_467_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_109_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311o_2 VPB VNB VGND VPWR C1 B1 A1 A2 A3 X
X0 a_79_21# C1 a_635_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.21 ps=1.42 w=1 l=0.15
X1 VPWR A2 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.17 ps=1.34 w=1 l=0.15
X2 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.13325 ps=1.06 w=0.65 l=0.15
X3 a_417_47# A2 a_319_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.1105 ps=0.99 w=0.65 l=0.15
X4 a_79_21# A1 a_417_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12025 ps=1.02 w=0.65 l=0.15
X5 a_319_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.156 ps=1.13 w=0.65 l=0.15
X6 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.24 pd=1.48 as=0.135 ps=1.27 w=1 l=0.15
X7 a_319_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.185 ps=1.37 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.156 pd=1.13 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_319_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.34 as=0.24 ps=1.48 w=1 l=0.15
X10 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13975 ps=1.08 w=0.65 l=0.15
X11 a_635_297# B1 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.21 ps=1.42 w=1 l=0.15
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_2 VPWR VGND VNB VPB A_N B C D X
X0 VPWR a_193_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# a_27_413# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.103975 ps=1 w=0.65 l=0.15
X4 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14325 pd=1.33 as=0.06615 ps=0.735 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103975 pd=1 as=0.06195 ps=0.715 w=0.42 l=0.15
X7 VGND a_193_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X8 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X9 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X10 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.14325 ps=1.33 w=1 l=0.15
X11 a_193_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0735 ps=0.77 w=0.42 l=0.15
X13 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4bb_2 VPWR VGND VPB VNB B A C_N D_N X
X0 a_398_413# a_206_93# a_316_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1215 pd=1.33 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VPWR a_316_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_316_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X3 X a_316_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X4 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1226 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND a_27_410# a_316_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X7 VGND A a_316_413# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND a_316_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_566_297# B a_494_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05985 pd=0.705 as=0.0441 ps=0.63 w=0.42 l=0.15
X10 a_206_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06195 ps=0.715 w=0.42 l=0.15
X11 a_316_413# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_206_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1226 ps=1.32 w=0.42 l=0.15
X13 a_494_297# a_27_410# a_398_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1215 ps=1.33 w=0.42 l=0.15
X14 a_316_413# a_206_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X15 VPWR A a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.05985 ps=0.705 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3b_2 VNB VPB VGND VPWR A_N C B Y
X0 a_408_47# B a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_408_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y a_27_47# a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17575 pd=1.395 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND C a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 a_218_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11975 ps=1.045 w=0.65 l=0.15
X7 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_218_47# B a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.17575 ps=1.395 w=1 l=0.15
X12 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11975 pd=1.045 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a41o_2 VNB VPB VGND VPWR X A1 A2 A3 A4 B1
X0 a_381_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A2 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X2 a_465_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_549_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13975 ps=1.08 w=0.65 l=0.15
X7 a_381_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A4 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_381_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 a_79_21# A1 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41a_2 VNB VPB VGND VPWR A1 A2 A3 A4 B1 X
X0 VGND A2 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.11375 ps=1 w=0.65 l=0.15
X1 a_496_297# A4 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.3025 ps=1.605 w=1 l=0.15
X2 a_393_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.115375 ps=1.005 w=0.65 l=0.15
X3 VPWR A1 a_697_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=2.82 as=0.175 ps=1.35 w=1 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3025 pd=1.605 as=0.305 ps=1.61 w=1 l=0.15
X7 VGND A4 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.118625 ps=1.015 w=0.65 l=0.15
X8 a_697_297# A2 a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X9 a_393_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2665 pd=2.12 as=0.11375 ps=1 w=0.65 l=0.15
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_393_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.208 ps=1.94 w=0.65 l=0.15
X12 a_597_297# A3 a_496_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.1775 ps=1.355 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_2 VNB VPB VGND VPWR A2 A1 B1_N X
X0 VGND B1_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND A2 a_478_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.105625 ps=0.975 w=0.65 l=0.15
X2 a_478_47# a_27_93# a_174_21# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_478_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X7 VPWR A1 a_574_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X8 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR B1_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 a_574_297# A2 a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X11 a_174_21# a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.395 ps=1.79 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_2 VNB VPB VGND VPWR A_N Y B
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X1 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.194 pd=1.95 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND B a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y a_27_93# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_229_47# a_27_93# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1468 ps=1.34 w=1 l=0.15
X6 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.165 ps=1.33 w=1 l=0.15
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X8 a_229_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1468 pd=1.34 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221oi_2 VNB VPB VGND VPWR A2 A1 B1 B2 Y C1
X0 Y B1 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_301_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_301_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND B2 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A1 a_735_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_297# B2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR A1 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_735_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_301_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1755 ps=1.84 w=0.65 l=0.15
X12 VPWR A2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X13 a_383_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X14 a_383_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_735_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X16 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X17 a_301_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X18 a_735_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B1 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_2 VPWR VGND VPB VNB A2 A1 Y B1 C1
X0 VGND A2 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR A1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_37_297# B1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_485_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_292_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VPWR A2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_485_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X11 a_37_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 Y A1 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X13 Y C1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14 a_292_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15 a_292_297# B1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_2 VPB VNB VGND VPWR A Y C_N B
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND a_531_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR C_N a_531_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9 a_281_297# a_531_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X10 Y a_531_21# a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 VGND C_N a_531_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X13 Y a_531_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111ai_2 VNB VPB VPWR VGND D1 Y C1 B1 A1 A2
X0 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_298_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VGND A1 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3 a_664_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND A2 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_298_47# B1 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.1755 ps=1.84 w=0.65 l=0.15
X7 a_497_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.22425 ps=1.99 w=0.65 l=0.15
X9 a_497_47# B1 a_298_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 Y A2 a_664_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.295 ps=2.59 w=1 l=0.15
X12 a_27_47# C1 a_298_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.091 ps=0.93 w=0.65 l=0.15
X13 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X16 a_497_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.091 ps=0.93 w=0.65 l=0.15
X17 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X18 VPWR A1 a_664_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 a_664_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_2 VNB VPB VPWR VGND B1_N A2 Y A1
X0 Y a_61_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183125 ps=1.24 w=0.65 l=0.15
X1 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_217_297# a_61_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_479_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 a_217_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5 Y a_61_47# a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR A1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_61_47# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X8 VGND A2 a_637_47# VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND a_61_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A1 a_479_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.06825 ps=0.86 w=0.65 l=0.15
X11 VGND B1_N a_61_47# VNB sky130_fd_pr__nfet_01v8 ad=0.183125 pd=1.24 as=0.126 ps=1.44 w=0.42 l=0.15
X12 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X13 a_637_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_2 VNB VPB VPWR VGND A_N X B
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.22895 ps=1.745 w=1 l=0.15
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22895 pd=1.745 as=0.0609 ps=0.71 w=0.42 l=0.15
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311ai_2 VGND VPWR VPB VNB Y B1 C1 A1 A2 A3
X0 VPWR A1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 a_55_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y C1 a_729_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.205 ps=1.41 w=1 l=0.15
X4 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_55_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.23075 ps=1.36 w=0.65 l=0.15
X6 VGND A1 a_55_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 a_55_47# B1 a_729_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND A2 a_55_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.305 ps=1.61 w=1 l=0.15
X10 VGND A3 a_55_47# VNB sky130_fd_pr__nfet_01v8 ad=0.23075 pd=1.36 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_729_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X12 a_51_297# A2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13 a_729_47# B1 a_55_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_301_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_55_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X17 a_51_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 Y A3 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_301_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4b_2 VNB VPB VGND VPWR A_N Y B C D
X0 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_465_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND D a_655_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X3 a_215_47# B a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_655_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_655_47# C a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.37 pd=1.74 as=0.135 ps=1.27 w=1 l=0.15
X8 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_465_47# C a_655_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=2.8 as=0.135 ps=1.27 w=1 l=0.15
X13 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.18 ps=1.36 w=1 l=0.15
X14 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.37 ps=1.74 w=1 l=0.15
X17 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111a_2 VPB VNB VGND VPWR X D1 C1 B1 A2 A1
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 a_80_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.365 ps=1.73 w=1 l=0.15
X3 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VPWR C1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.14 ps=1.28 w=1 l=0.15
X5 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X6 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X7 a_674_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X8 a_386_47# D1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X9 VPWR A1 a_674_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.195 ps=1.39 w=1 l=0.15
X10 a_566_47# B1 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X11 VGND A2 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X12 a_566_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X13 a_458_47# C1 a_386_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
.ends

.subckt aes_core VGND VPWR block[0] block[100] block[101] block[102] block[103] block[104]
+ block[105] block[106] block[107] block[108] block[109] block[10] block[110] block[111]
+ block[112] block[113] block[114] block[115] block[116] block[117] block[118] block[119]
+ block[11] block[120] block[121] block[122] block[123] block[124] block[125] block[126]
+ block[127] block[12] block[13] block[14] block[15] block[16] block[17] block[18]
+ block[19] block[1] block[20] block[21] block[22] block[23] block[24] block[25] block[26]
+ block[27] block[28] block[29] block[2] block[30] block[31] block[32] block[33] block[34]
+ block[35] block[36] block[37] block[38] block[39] block[3] block[40] block[41] block[42]
+ block[43] block[44] block[45] block[46] block[47] block[48] block[49] block[4] block[50]
+ block[51] block[52] block[53] block[54] block[55] block[56] block[57] block[58]
+ block[59] block[5] block[60] block[61] block[62] block[63] block[64] block[65] block[66]
+ block[67] block[68] block[69] block[6] block[70] block[71] block[72] block[73] block[74]
+ block[75] block[76] block[77] block[78] block[79] block[7] block[80] block[81] block[82]
+ block[83] block[84] block[85] block[86] block[87] block[88] block[89] block[8] block[90]
+ block[91] block[92] block[93] block[94] block[95] block[96] block[97] block[98]
+ block[99] block[9] clk encdec init key[0] key[100] key[101] key[102] key[103] key[104]
+ key[105] key[106] key[107] key[108] key[109] key[10] key[110] key[111] key[112]
+ key[113] key[114] key[115] key[116] key[117] key[118] key[119] key[11] key[120]
+ key[121] key[122] key[123] key[124] key[125] key[126] key[127] key[128] key[129]
+ key[12] key[130] key[131] key[132] key[133] key[134] key[135] key[136] key[137]
+ key[138] key[139] key[13] key[140] key[141] key[142] key[143] key[144] key[145]
+ key[146] key[147] key[148] key[149] key[14] key[150] key[151] key[152] key[153]
+ key[154] key[155] key[156] key[157] key[158] key[159] key[15] key[160] key[161]
+ key[162] key[163] key[164] key[165] key[166] key[167] key[168] key[169] key[16]
+ key[170] key[171] key[172] key[173] key[174] key[175] key[176] key[177] key[178]
+ key[179] key[17] key[180] key[181] key[182] key[183] key[184] key[185] key[186]
+ key[187] key[188] key[189] key[18] key[190] key[191] key[192] key[193] key[194]
+ key[195] key[196] key[197] key[198] key[199] key[19] key[1] key[200] key[201] key[202]
+ key[203] key[204] key[205] key[206] key[207] key[208] key[209] key[20] key[210]
+ key[211] key[212] key[213] key[214] key[215] key[216] key[217] key[218] key[219]
+ key[21] key[220] key[221] key[222] key[223] key[224] key[225] key[226] key[227]
+ key[228] key[229] key[22] key[230] key[231] key[232] key[233] key[234] key[235]
+ key[236] key[237] key[238] key[239] key[23] key[240] key[241] key[242] key[243]
+ key[244] key[245] key[246] key[247] key[248] key[249] key[24] key[250] key[251]
+ key[252] key[253] key[254] key[255] key[25] key[26] key[27] key[28] key[29] key[2]
+ key[30] key[31] key[32] key[33] key[34] key[35] key[36] key[37] key[38] key[39]
+ key[3] key[40] key[41] key[42] key[43] key[44] key[45] key[46] key[47] key[48] key[49]
+ key[4] key[50] key[51] key[52] key[53] key[54] key[55] key[56] key[57] key[58] key[59]
+ key[5] key[60] key[61] key[62] key[63] key[64] key[65] key[66] key[67] key[68] key[69]
+ key[6] key[70] key[71] key[72] key[73] key[74] key[75] key[76] key[77] key[78] key[79]
+ key[7] key[80] key[81] key[82] key[83] key[84] key[85] key[86] key[87] key[88] key[89]
+ key[8] key[90] key[91] key[92] key[93] key[94] key[95] key[96] key[97] key[98] key[99]
+ key[9] keylen next ready reset_n result[0] result[100] result[101] result[102] result[103]
+ result[104] result[105] result[106] result[107] result[108] result[109] result[10]
+ result[110] result[111] result[112] result[113] result[114] result[115] result[116]
+ result[117] result[118] result[119] result[11] result[120] result[121] result[122]
+ result[123] result[124] result[125] result[126] result[127] result[12] result[13]
+ result[14] result[15] result[16] result[17] result[18] result[19] result[1] result[20]
+ result[21] result[22] result[23] result[24] result[25] result[26] result[27] result[28]
+ result[29] result[2] result[30] result[31] result[32] result[33] result[34] result[35]
+ result[36] result[37] result[38] result[39] result[3] result[40] result[41] result[42]
+ result[43] result[44] result[45] result[46] result[47] result[48] result[49] result[4]
+ result[50] result[51] result[52] result[53] result[54] result[55] result[56] result[57]
+ result[58] result[59] result[5] result[60] result[61] result[62] result[63] result[64]
+ result[65] result[66] result[67] result[68] result[69] result[6] result[70] result[71]
+ result[72] result[73] result[74] result[75] result[76] result[77] result[78] result[79]
+ result[7] result[80] result[81] result[82] result[83] result[84] result[85] result[86]
+ result[87] result[88] result[89] result[8] result[90] result[91] result[92] result[93]
+ result[94] result[95] result[96] result[97] result[98] result[99] result[9] result_valid
XFILLER_0_158_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_253_367 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18869_ VGND VPWR _04713_ _04710_ _04712_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20900_ VGND VPWR VGND VPWR _05895_ keymem.key_mem_we _03150_ _05893_ _01200_ sky130_fd_sc_hd__a31o_2
XFILLER_0_27_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21880_ VPWR VGND keymem.key_mem\[3\]\[8\] _06416_ _06413_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_136_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20831_ VGND VPWR VGND VPWR _05858_ keymem.key_mem_we _02787_ _05850_ _01168_ sky130_fd_sc_hd__a31o_2
XFILLER_0_72_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23550_ VGND VPWR VPWR VGND clk _00051_ reset_n keymem.key_mem\[14\]\[39\] sky130_fd_sc_hd__dfrtp_2
X_20762_ VPWR VGND VGND VPWR _05818_ keymem.round_ctr_reg\[2\] _05241_ sky130_fd_sc_hd__nand2_2
XFILLER_0_33_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1342 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_159_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22501_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[50\] _06737_ _06736_ _04955_ _01958_
+ sky130_fd_sc_hd__a22o_2
X_23481_ VGND VPWR _07343_ enc_block.block_w0_reg\[21\] _07283_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20693_ VGND VPWR VPWR VGND _05772_ _03459_ keymem.key_mem\[8\]\[95\] _05782_ sky130_fd_sc_hd__mux2_2
X_25220_ VGND VPWR VPWR VGND clk _01713_ reset_n keymem.key_mem\[3\]\[61\] sky130_fd_sc_hd__dfrtp_2
X_22432_ VGND VPWR VPWR VGND _06702_ keymem.key_mem\[1\]\[10\] _10836_ _06710_ sky130_fd_sc_hd__mux2_2
XFILLER_0_9_499 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_169_1263 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_247_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25151_ VGND VPWR VPWR VGND clk _01644_ reset_n keymem.key_mem\[4\]\[120\] sky130_fd_sc_hd__dfrtp_2
X_22363_ VGND VPWR _01886_ _06672_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_245_1151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24102_ VGND VPWR VPWR VGND clk _00595_ reset_n keymem.key_mem\[12\]\[95\] sky130_fd_sc_hd__dfrtp_2
X_21314_ VGND VPWR _06114_ _06113_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_143_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25082_ VGND VPWR VPWR VGND clk _01575_ reset_n keymem.key_mem\[4\]\[51\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_694 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22294_ VGND VPWR _01853_ _06636_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_182_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_973 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_770 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_83_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24033_ VGND VPWR VPWR VGND clk _00526_ reset_n keymem.key_mem\[12\]\[26\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_143_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21245_ VGND VPWR VPWR VGND _06076_ _03459_ keymem.key_mem\[6\]\[95\] _06078_ sky130_fd_sc_hd__mux2_2
XFILLER_0_13_483 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_110_2_Left_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21176_ VGND VPWR VPWR VGND _06040_ _03172_ keymem.key_mem\[6\]\[62\] _06042_ sky130_fd_sc_hd__mux2_2
XFILLER_0_223_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20127_ VGND VPWR VPWR VGND _05482_ _03364_ keymem.key_mem\[10\]\[84\] _05483_ sky130_fd_sc_hd__mux2_2
XFILLER_0_256_183 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_245_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20058_ VGND VPWR VPWR VGND _05446_ _03068_ keymem.key_mem\[10\]\[51\] _05447_ sky130_fd_sc_hd__mux2_2
X_24935_ VGND VPWR VPWR VGND clk _01428_ reset_n keymem.key_mem\[5\]\[32\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_176_1256 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_99_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_242_Right_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11900_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[21\] dec_new_block\[117\]
+ _07514_ sky130_fd_sc_hd__mux2_2
X_24866_ VGND VPWR VPWR VGND clk _01359_ reset_n keymem.key_mem\[6\]\[91\] sky130_fd_sc_hd__dfrtp_2
X_12880_ VGND VPWR VGND VPWR _08412_ _08050_ keymem.key_mem\[7\]\[71\] _08409_ _08411_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_217_1242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_161_1_Left_428 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_154_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11831_ VGND VPWR result[82] _07479_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23817_ VGND VPWR VPWR VGND clk _00310_ reset_n enc_block.block_w1_reg\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_90_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_150_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24797_ VGND VPWR VPWR VGND clk _01290_ reset_n keymem.key_mem\[6\]\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_261_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1061 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14550_ VPWR VGND VPWR VGND _10013_ _10017_ _10015_ _09195_ _10018_ sky130_fd_sc_hd__or4_2
XFILLER_0_90_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11762_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[16\] dec_new_block\[48\]
+ _07445_ sky130_fd_sc_hd__mux2_2
X_23748_ keymem.prev_key0_reg\[104\] clk _00245_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_51_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13501_ VPWR VGND VGND VPWR enc_block.block_w1_reg\[7\] enc_block.sword_ctr_reg\[0\]
+ _08973_ sky130_fd_sc_hd__or2b_2
XFILLER_0_55_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14481_ VGND VPWR VGND VPWR _09089_ _09137_ _09124_ _09115_ _09950_ sky130_fd_sc_hd__o22a_2
X_23679_ keymem.prev_key0_reg\[35\] clk _00176_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_11693_ VGND VPWR result[13] _07410_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_265_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_230_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16220_ VPWR VGND VGND VPWR _11361_ _02385_ _11252_ sky130_fd_sc_hd__nor2_2
X_13432_ VPWR VGND VPWR VGND _08908_ keymem.key_mem\[14\]\[126\] _07963_ keymem.key_mem\[6\]\[126\]
+ _08137_ _08909_ sky130_fd_sc_hd__a221o_2
X_25418_ VGND VPWR VPWR VGND clk _01911_ reset_n keymem.key_mem\[1\]\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_187_1352 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16151_ VGND VPWR VGND VPWR _11278_ _11604_ _11250_ _11469_ _11605_ sky130_fd_sc_hd__o22a_2
XFILLER_0_118_290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25349_ VGND VPWR VPWR VGND clk _01842_ reset_n keymem.key_mem\[2\]\[62\] sky130_fd_sc_hd__dfrtp_2
X_13363_ VGND VPWR VGND VPWR _08847_ _07912_ keymem.key_mem\[11\]\[119\] _08844_ _08846_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_23_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15102_ VGND VPWR _10566_ _10540_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_51_556 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12314_ VPWR VGND VPWR VGND keymem.key_mem\[4\]\[19\] _07854_ keymem.key_mem\[2\]\[19\]
+ _07647_ _07898_ sky130_fd_sc_hd__a22o_2
XFILLER_0_161_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16082_ VGND VPWR _11537_ keymem.prev_key0_reg\[49\] keymem.prev_key0_reg\[81\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_263_1273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13294_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[112\] _08714_ _08784_ _08780_ _08785_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_133_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_415 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_210_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15033_ VPWR VGND VPWR VGND _10473_ _10477_ _10453_ _10451_ _10497_ sky130_fd_sc_hd__or4_2
XFILLER_0_224_1257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19910_ VGND VPWR VPWR VGND _05361_ keymem.key_mem\[11\]\[111\] _03560_ _05367_ sky130_fd_sc_hd__mux2_2
XFILLER_0_161_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12245_ VGND VPWR _07834_ _07694_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_48_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19841_ VGND VPWR VPWR VGND _05328_ keymem.key_mem\[11\]\[78\] _03314_ _05331_ sky130_fd_sc_hd__mux2_2
XFILLER_0_202_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12176_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[9\] _07609_ keymem.key_mem\[10\]\[9\]
+ _07561_ _07770_ sky130_fd_sc_hd__a22o_2
XFILLER_0_202_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19772_ VGND VPWR VPWR VGND _05292_ keymem.key_mem\[11\]\[45\] _03006_ _05295_ sky130_fd_sc_hd__mux2_2
X_16984_ VPWR VGND _03111_ _02703_ _02702_ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_263_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15935_ VPWR VGND VGND VPWR _11391_ _11180_ _11258_ sky130_fd_sc_hd__nand2_2
X_18723_ VPWR VGND VPWR VGND _04580_ block[94] _04576_ enc_block.block_w1_reg\[30\]
+ _04543_ _04581_ sky130_fd_sc_hd__a221o_2
XFILLER_0_155_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18654_ VPWR VGND _04520_ _04519_ enc_block.round_key\[86\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15866_ VGND VPWR VGND VPWR _11321_ _11315_ _11322_ _11310_ _11309_ sky130_fd_sc_hd__nand4_2
XFILLER_0_64_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_612 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14817_ VPWR VGND VPWR VGND _10282_ _10085_ _10271_ key[134] _09544_ _10283_ sky130_fd_sc_hd__a221o_2
X_17605_ VGND VPWR _00138_ _03662_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18585_ VPWR VGND _04458_ _04457_ enc_block.round_key\[79\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15797_ VGND VPWR _11253_ _11252_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_15_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17536_ VGND VPWR VPWR VGND _02588_ _02589_ _09932_ _03602_ sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_186_2_Left_657 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_147_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14748_ VGND VPWR VGND VPWR _09640_ _09704_ _10211_ _10214_ _10213_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_50_1003 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_15_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_58_188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17467_ VPWR VGND VPWR VGND _03542_ _03494_ _03540_ key[236] _03527_ _03543_ sky130_fd_sc_hd__a221o_2
XFILLER_0_11_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14679_ VGND VPWR _10146_ keymem.prev_key0_reg\[37\] keymem.prev_key0_reg\[69\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_156_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_89_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16418_ VPWR VGND VGND VPWR _11222_ _11203_ _02580_ _11325_ _11370_ _11275_ sky130_fd_sc_hd__o32ai_2
XFILLER_0_251_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19206_ VPWR VGND keymem.key_mem\[13\]\[60\] _04970_ _04961_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_73_158 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17398_ VGND VPWR VPWR VGND _09730_ _09925_ key[227] _03483_ sky130_fd_sc_hd__mux2_2
XFILLER_0_89_1279 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_116_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19137_ VPWR VGND keymem.key_mem\[13\]\[35\] _04926_ _04915_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16349_ VGND VPWR VGND VPWR _11298_ _11302_ _11361_ _11344_ _02512_ sky130_fd_sc_hd__o22a_2
XFILLER_0_89_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_42_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_1_Right_676 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19068_ VGND VPWR VGND VPWR _04886_ keymem.key_mem_we _10194_ _04878_ _00377_ sky130_fd_sc_hd__a31o_2
XFILLER_0_120_63 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_129_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_120_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18019_ VGND VPWR VGND VPWR _03941_ enc_block.round\[1\] _03944_ enc_block.round\[2\]
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_242_1357 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_22_280 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21030_ VGND VPWR _01262_ _05963_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_22_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_971 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_125_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_196_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1081 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_22_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_96_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22981_ VGND VPWR _02996_ _02990_ _06956_ _02991_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_198_219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_59_1061 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24720_ VGND VPWR VPWR VGND clk _01213_ reset_n keymem.key_mem\[7\]\[73\] sky130_fd_sc_hd__dfrtp_2
X_21932_ VGND VPWR VPWR VGND _06403_ _04920_ keymem.key_mem\[3\]\[32\] _06444_ sky130_fd_sc_hd__mux2_2
XFILLER_0_59_1083 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24651_ VGND VPWR VPWR VGND clk _01144_ reset_n keymem.key_mem\[7\]\[4\] sky130_fd_sc_hd__dfrtp_2
X_21863_ VPWR VGND keymem.key_mem\[3\]\[0\] _06407_ _06406_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_33_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23602_ VGND VPWR VPWR VGND clk _00103_ reset_n keymem.key_mem\[14\]\[91\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_136_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20814_ VPWR VGND keymem.key_mem\[7\]\[21\] _05849_ _05844_ VPWR VGND sky130_fd_sc_hd__and2_2
X_24582_ VGND VPWR VPWR VGND clk _01075_ reset_n keymem.key_mem\[8\]\[63\] sky130_fd_sc_hd__dfrtp_2
X_21794_ VGND VPWR _01621_ _06368_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_72_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23533_ VGND VPWR VPWR VGND clk _00034_ reset_n keymem.key_mem\[14\]\[22\] sky130_fd_sc_hd__dfrtp_2
X_20745_ VGND VPWR _01131_ _05809_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_212_1172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_18_553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23464_ VGND VPWR _07328_ _07274_ _07327_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_68_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20676_ VGND VPWR _01098_ _05773_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_64_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_174_182 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_107_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25203_ VGND VPWR VPWR VGND clk _01696_ reset_n keymem.key_mem\[3\]\[44\] sky130_fd_sc_hd__dfrtp_2
X_22415_ VGND VPWR VPWR VGND _06696_ keymem.key_mem\[1\]\[3\] _09992_ _06700_ sky130_fd_sc_hd__mux2_2
X_23395_ VGND VPWR _07267_ enc_block.block_w0_reg\[23\] _07266_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25134_ VGND VPWR VPWR VGND clk _01627_ reset_n keymem.key_mem\[4\]\[103\] sky130_fd_sc_hd__dfrtp_2
X_22346_ VGND VPWR _01878_ _06663_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_108_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_143_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22277_ VGND VPWR _01845_ _06627_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25065_ VGND VPWR VPWR VGND clk _01558_ reset_n keymem.key_mem\[4\]\[34\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_108_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12030_ VGND VPWR _07631_ _07599_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21228_ VGND VPWR VPWR VGND _06065_ _03392_ keymem.key_mem\[6\]\[87\] _06069_ sky130_fd_sc_hd__mux2_2
X_24016_ VGND VPWR VPWR VGND clk _00509_ reset_n keymem.key_mem\[12\]\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_104_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_835 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21159_ VGND VPWR VPWR VGND _06029_ _03090_ keymem.key_mem\[6\]\[54\] _06033_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_665 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_79_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13981_ VPWR VGND VGND VPWR _09452_ _09453_ _09355_ sky130_fd_sc_hd__nor2_2
XFILLER_0_254_1217 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_217_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_258_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15720_ VGND VPWR VGND VPWR _11176_ enc_block.sword_ctr_reg\[0\] enc_block.block_w1_reg\[17\]
+ enc_block.sword_ctr_reg\[1\] sky130_fd_sc_hd__and3b_2
XFILLER_0_244_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12932_ VGND VPWR enc_block.round_key\[76\] _08458_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24918_ VGND VPWR VPWR VGND clk _01411_ reset_n keymem.key_mem\[5\]\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_125_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15651_ VGND VPWR VPWR VGND _11107_ _11103_ _11102_ _11108_ sky130_fd_sc_hd__mux2_2
XFILLER_0_119_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_154_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12863_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[70\] _08137_ keymem.key_mem\[2\]\[70\]
+ _08116_ _08396_ sky130_fd_sc_hd__a22o_2
X_24849_ VGND VPWR VPWR VGND clk _01342_ reset_n keymem.key_mem\[6\]\[74\] sky130_fd_sc_hd__dfrtp_2
X_14602_ VGND VPWR VPWR VGND _09751_ _10069_ _09747_ _10070_ sky130_fd_sc_hd__or3_2
XFILLER_0_115_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18370_ VGND VPWR _04265_ enc_block.round_key\[123\] _04264_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_11814_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[10\] dec_new_block\[74\]
+ _07471_ sky130_fd_sc_hd__mux2_2
XFILLER_0_154_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15582_ VGND VPWR _11041_ _09863_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_95_250 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12794_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[63\] _07812_ keymem.key_mem\[12\]\[63\]
+ _07806_ _08334_ sky130_fd_sc_hd__a22o_2
XFILLER_0_51_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_626 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_115_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17321_ VPWR VGND VPWR VGND _03415_ key[90] _11543_ sky130_fd_sc_hd__or2_2
XFILLER_0_16_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14533_ VGND VPWR VGND VPWR _09054_ _09181_ _09998_ _09999_ _10001_ _10000_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_189_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11745_ VGND VPWR result[39] _07436_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_230_1261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17252_ VGND VPWR _03352_ _10967_ _03353_ _02403_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_55_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14464_ VGND VPWR _09933_ keymem.prev_key0_reg\[35\] keymem.prev_key0_reg\[67\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_153_311 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_55_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_86_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11676_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[5\] dec_new_block\[5\]
+ _07402_ sky130_fd_sc_hd__mux2_2
XFILLER_0_165_182 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16203_ VPWR VGND VPWR VGND _02365_ _02367_ _02366_ _02364_ _02368_ sky130_fd_sc_hd__or4_2
XFILLER_0_187_1171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_372 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13415_ VGND VPWR enc_block.round_key\[124\] _08893_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_265_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17183_ VGND VPWR VPWR VGND _02864_ _10963_ keymem.prev_key0_reg\[76\] _03291_ sky130_fd_sc_hd__or3_2
X_14395_ VGND VPWR VPWR VGND _09864_ keymem.key_mem\[14\]\[2\] _09862_ _09865_ sky130_fd_sc_hd__mux2_2
XFILLER_0_3_417 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16134_ VGND VPWR VPWR VGND _11306_ _11464_ _11588_ _11587_ _11584_ sky130_fd_sc_hd__o211a_2
XFILLER_0_24_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1010 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13346_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[118\] _08009_ keymem.key_mem\[11\]\[118\]
+ _08011_ _08831_ sky130_fd_sc_hd__a22o_2
XFILLER_0_24_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_126_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16065_ VGND VPWR VGND VPWR _11276_ _11412_ _11512_ _11515_ _11520_ _11519_ sky130_fd_sc_hd__a2111o_2
X_13277_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[111\] _07703_ keymem.key_mem\[12\]\[111\]
+ _07788_ _08769_ sky130_fd_sc_hd__a22o_2
XFILLER_0_59_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_126_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15016_ VGND VPWR _10480_ _10437_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_122_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12228_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[12\] _07568_ keymem.key_mem\[14\]\[12\]
+ _07632_ _07819_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_835 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_166_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19824_ VGND VPWR VPWR VGND _05314_ keymem.key_mem\[11\]\[70\] _03245_ _05322_ sky130_fd_sc_hd__mux2_2
XFILLER_0_23_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12159_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[8\] _07619_ keymem.key_mem\[8\]\[8\]
+ _07753_ _07754_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_118_2_Right_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_209_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19755_ VGND VPWR VPWR VGND _05281_ keymem.key_mem\[11\]\[37\] _02924_ _05286_ sky130_fd_sc_hd__mux2_2
X_16967_ VGND VPWR VPWR VGND _09511_ key[183] keymem.prev_key1_reg\[55\] _03096_ sky130_fd_sc_hd__mux2_2
XFILLER_0_237_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_890 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18706_ VPWR VGND VPWR VGND _04565_ block[92] _04487_ enc_block.block_w1_reg\[28\]
+ _04543_ _04566_ sky130_fd_sc_hd__a221o_2
XFILLER_0_264_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15918_ VPWR VGND VPWR VGND _11371_ _11373_ _11374_ _11366_ _11368_ sky130_fd_sc_hd__or4b_2
XFILLER_0_56_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19686_ VGND VPWR VPWR VGND _05247_ keymem.key_mem\[11\]\[4\] _10099_ _05250_ sky130_fd_sc_hd__mux2_2
X_16898_ VGND VPWR VGND VPWR keylen _03034_ _03033_ keymem.prev_key1_reg\[48\] _11154_
+ _11155_ sky130_fd_sc_hd__a311oi_2
X_15849_ VGND VPWR _11305_ _11304_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18637_ VGND VPWR _04504_ _03952_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_172_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_133_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18568_ VGND VPWR VGND VPWR _04441_ _03951_ _04442_ _00321_ sky130_fd_sc_hd__a21o_2
XFILLER_0_34_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_272 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17519_ VPWR VGND VGND VPWR _03587_ _02460_ _02461_ sky130_fd_sc_hd__nand2_2
X_18499_ VPWR VGND VGND VPWR _04380_ _04381_ _04052_ sky130_fd_sc_hd__nor2_2
XFILLER_0_213_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20530_ VGND VPWR VPWR VGND _05692_ _11546_ keymem.key_mem\[8\]\[17\] _05697_ sky130_fd_sc_hd__mux2_2
XFILLER_0_28_862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20461_ VGND VPWR _00997_ _05659_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_248_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_54_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22200_ VGND VPWR VPWR VGND _06578_ _02811_ keymem.key_mem\[2\]\[29\] _06587_ sky130_fd_sc_hd__mux2_2
X_23180_ VGND VPWR VPWR VGND _02299_ _03630_ _03632_ _06976_ _07076_ sky130_fd_sc_hd__o31a_2
X_20392_ VGND VPWR _00964_ _05623_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_259_724 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_144_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22131_ VGND VPWR VPWR VGND _06402_ _05087_ keymem.key_mem\[3\]\[126\] _06549_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_76_1_Right_677 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_105_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22062_ VPWR VGND keymem.key_mem\[3\]\[93\] _06513_ _06405_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_80_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21013_ VGND VPWR _01254_ _05954_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_41_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25821_ VGND VPWR VPWR VGND clk _02314_ reset_n enc_block.block_w3_reg\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_255_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_890 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25752_ keymem.prev_key1_reg\[68\] clk _02245_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22964_ VGND VPWR _02922_ keylen _06946_ _02917_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_74_1334 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24703_ VGND VPWR VPWR VGND clk _01196_ reset_n keymem.key_mem\[7\]\[56\] sky130_fd_sc_hd__dfrtp_2
X_21915_ VPWR VGND keymem.key_mem\[3\]\[24\] _06435_ _06427_ VPWR VGND sky130_fd_sc_hd__and2_2
X_25683_ VGND VPWR VPWR VGND clk _02176_ reset_n keymem.ready sky130_fd_sc_hd__dfrtp_2
X_22895_ VGND VPWR VGND VPWR _06903_ _10901_ _06891_ _10912_ _06892_ sky130_fd_sc_hd__a211o_2
XFILLER_0_253_1272 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24634_ VGND VPWR VPWR VGND clk _01127_ reset_n keymem.key_mem\[8\]\[115\] sky130_fd_sc_hd__dfrtp_2
X_21846_ VGND VPWR _01646_ _06395_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_77_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24565_ VGND VPWR VPWR VGND clk _01058_ reset_n keymem.key_mem\[8\]\[46\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_231_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21777_ VGND VPWR _01613_ _06359_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_4_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23516_ VGND VPWR VPWR VGND clk _00017_ reset_n keymem.key_mem\[14\]\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_862 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_92_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20728_ VGND VPWR _01123_ _05800_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_4_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24496_ VGND VPWR VPWR VGND clk _00989_ reset_n keymem.key_mem\[9\]\[105\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_147_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_92_286 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_162_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23447_ VPWR VGND VGND VPWR _07313_ _07247_ _07312_ sky130_fd_sc_hd__nand2_2
X_20659_ VGND VPWR _01090_ _05764_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_34_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1076 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13200_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[103\] _07622_ keymem.key_mem\[4\]\[103\]
+ _07637_ _08700_ sky130_fd_sc_hd__a22o_2
X_14180_ VPWR VGND VGND VPWR _09082_ _09651_ _09033_ sky130_fd_sc_hd__nor2_2
X_23378_ _07250_ _07252_ _04103_ _07251_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_33_375 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25117_ VGND VPWR VPWR VGND clk _01610_ reset_n keymem.key_mem\[4\]\[86\] sky130_fd_sc_hd__dfrtp_2
X_13131_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[96\] _07583_ keymem.key_mem\[6\]\[96\]
+ _07771_ _08638_ sky130_fd_sc_hd__a22o_2
X_22329_ VGND VPWR _01870_ _06654_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_108_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13062_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[89\] _08449_ _08575_ _08571_ _08576_
+ sky130_fd_sc_hd__o22a_2
X_25048_ VGND VPWR VPWR VGND clk _01541_ reset_n keymem.key_mem\[4\]\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_29_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12013_ VPWR VGND VPWR VGND _07614_ keymem.key_mem\[5\]\[1\] _07613_ keymem.key_mem\[9\]\[1\]
+ _07612_ _07615_ sky130_fd_sc_hd__a221o_2
X_17870_ VGND VPWR _00222_ _03843_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_264_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_79_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_105_1_Left_372 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_206_805 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16821_ VPWR VGND VPWR VGND _02963_ _02960_ _02958_ key[169] _02875_ _02964_ sky130_fd_sc_hd__a221o_2
XFILLER_0_79_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16752_ VGND VPWR VPWR VGND _02901_ _09985_ _09933_ _10735_ _02900_ sky130_fd_sc_hd__o31ai_2
X_19540_ VGND VPWR VPWR VGND _05151_ _04975_ keymem.key_mem\[12\]\[65\] _05171_ sky130_fd_sc_hd__mux2_2
X_13964_ _09364_ _09436_ _09332_ _09389_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_215_1009 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_214_860 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_232_167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_219_1189 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15703_ _11155_ _11159_ _11154_ _11156_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_12915_ VGND VPWR VGND VPWR _07912_ keymem.key_mem\[11\]\[75\] _08440_ _08442_ _08443_
+ _08243_ sky130_fd_sc_hd__a2111o_2
X_19471_ VGND VPWR VPWR VGND _05092_ _04922_ keymem.key_mem\[12\]\[33\] _05134_ sky130_fd_sc_hd__mux2_2
X_16683_ VPWR VGND VPWR VGND _02837_ _10325_ _02834_ _02835_ _02836_ _10281_ sky130_fd_sc_hd__o311a_2
X_13895_ VPWR VGND VGND VPWR _09366_ _09367_ _09268_ sky130_fd_sc_hd__nor2_2
XFILLER_0_213_370 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18422_ VPWR VGND VGND VPWR _04309_ _04310_ _03966_ sky130_fd_sc_hd__nor2_2
X_15634_ VGND VPWR _11092_ keymem.prev_key0_reg\[110\] _11091_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12846_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[68\] _07629_ keymem.key_mem\[1\]\[68\]
+ _07800_ _08381_ sky130_fd_sc_hd__a22o_2
XFILLER_0_57_913 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18353_ VPWR VGND VPWR VGND _04249_ _04189_ _04247_ enc_block.block_w0_reg\[25\]
+ _03993_ _00299_ sky130_fd_sc_hd__a221o_2
X_15565_ VGND VPWR VGND VPWR _11023_ _11021_ _11024_ _11022_ sky130_fd_sc_hd__nand3_2
XFILLER_0_185_266 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_16_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12777_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[61\] _07587_ keymem.key_mem\[11\]\[61\]
+ _07600_ _08319_ sky130_fd_sc_hd__a22o_2
X_17304_ VGND VPWR VGND VPWR keylen _03400_ _03399_ _10323_ _02681_ _02682_ sky130_fd_sc_hd__a311oi_2
X_14516_ VGND VPWR _09985_ keymem.prev_key0_reg\[99\] _09984_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_18284_ VPWR VGND VPWR VGND _04186_ block[115] _04076_ enc_block.block_w1_reg\[19\]
+ _04171_ _04187_ sky130_fd_sc_hd__a221o_2
X_11728_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[31\] dec_new_block\[31\]
+ _07428_ sky130_fd_sc_hd__mux2_2
X_15496_ VGND VPWR _10955_ _10527_ _10956_ _10867_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_9_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17235_ VGND VPWR VGND VPWR _03337_ _03042_ _03338_ keylen sky130_fd_sc_hd__a21oi_2
XFILLER_0_83_286 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14447_ VGND VPWR VGND VPWR _09452_ _09268_ _09916_ _09349_ sky130_fd_sc_hd__a21oi_2
X_11659_ VPWR VGND VPWR VGND _07393_ _07380_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_314 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_342 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17166_ VGND VPWR VGND VPWR _03275_ keylen _03273_ _03276_ _10902_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_25_887 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14378_ VGND VPWR VGND VPWR _09174_ _09136_ _09107_ _09019_ _09848_ sky130_fd_sc_hd__o22a_2
XFILLER_0_10_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16117_ VGND VPWR VGND VPWR _11296_ _11527_ _11473_ _11420_ _11571_ sky130_fd_sc_hd__o22a_2
X_13329_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[116\] _07649_ keymem.key_mem\[1\]\[116\]
+ _07714_ _08816_ sky130_fd_sc_hd__a22o_2
X_17097_ VGND VPWR VGND VPWR _03214_ _09513_ _10732_ key[67] sky130_fd_sc_hd__o21a_2
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_879 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16048_ VPWR VGND VGND VPWR _11275_ _11503_ _11396_ sky130_fd_sc_hd__nor2_2
XFILLER_0_126_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1226 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_97_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_900 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19807_ VGND VPWR VPWR VGND _05303_ keymem.key_mem\[11\]\[62\] _03173_ _05313_ sky130_fd_sc_hd__mux2_2
XFILLER_0_97_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_119_2_Right_191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17999_ VGND VPWR VGND VPWR _03737_ keymem.prev_key1_reg\[123\] _03931_ _03738_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_58_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19738_ VGND VPWR VPWR VGND _05270_ keymem.key_mem\[11\]\[29\] _02812_ _05277_ sky130_fd_sc_hd__mux2_2
XFILLER_0_223_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19669_ VGND VPWR _00626_ _05238_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21700_ VGND VPWR _06319_ _06262_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_35_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1086 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22680_ VGND VPWR VPWR VGND _06809_ keymem.key_mem\[0\]\[28\] _02787_ _06812_ sky130_fd_sc_hd__mux2_2
XFILLER_0_47_401 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21631_ VGND VPWR VPWR VGND _06275_ _02479_ keymem.key_mem\[4\]\[20\] _06283_ sky130_fd_sc_hd__mux2_2
XFILLER_0_34_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_168_1306 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_69_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24350_ VGND VPWR VPWR VGND clk _00843_ reset_n keymem.key_mem\[10\]\[87\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_191_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21562_ VGND VPWR _01512_ _06245_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_168_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_990 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23301_ VGND VPWR VGND VPWR _07182_ _04266_ _07095_ _07183_ enc_block.block_w3_reg\[9\]
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_69_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20513_ VGND VPWR VPWR VGND _05680_ _10746_ keymem.key_mem\[8\]\[9\] _05688_ sky130_fd_sc_hd__mux2_2
X_21493_ VGND VPWR _06209_ _06115_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24281_ VGND VPWR VPWR VGND clk _00774_ reset_n keymem.key_mem\[10\]\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_117_388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23232_ VGND VPWR _07120_ _07118_ _07119_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20444_ VGND VPWR VPWR VGND _05649_ _03525_ keymem.key_mem\[9\]\[105\] _05651_ sky130_fd_sc_hd__mux2_2
XFILLER_0_28_1111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_43_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23163_ VGND VPWR _02292_ _07066_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20375_ VGND VPWR VPWR VGND _05614_ _03259_ keymem.key_mem\[9\]\[72\] _05615_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_170_1_Left_437 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_105_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_1_Right_678 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22114_ VGND VPWR _01769_ _06540_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23094_ VGND VPWR VPWR VGND _06992_ _07022_ keymem.prev_key1_reg\[90\] _07023_ sky130_fd_sc_hd__mux2_2
XFILLER_0_100_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22045_ VGND VPWR _01736_ _06504_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_179_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_760 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_473 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_179_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25804_ keymem.prev_key1_reg\[120\] clk _02297_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_23996_ VGND VPWR VPWR VGND clk _00489_ reset_n keymem.key_mem\[13\]\[117\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_203_819 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_214_167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25735_ keymem.prev_key1_reg\[51\] clk _02228_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_253_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22947_ VGND VPWR VGND VPWR _02207_ _06935_ _06916_ keymem.prev_key1_reg\[30\] sky130_fd_sc_hd__o21a_2
XFILLER_0_74_1164 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12700_ VGND VPWR enc_block.round_key\[53\] _08249_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13680_ VPWR VGND VGND VPWR _09150_ _09041_ _09149_ _09146_ _09152_ _09151_ sky130_fd_sc_hd__o221a_2
X_25666_ VGND VPWR VPWR VGND clk _02159_ reset_n keymem.key_mem\[0\]\[123\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_116_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22878_ VGND VPWR VGND VPWR _06893_ _10084_ _06891_ _10097_ _06892_ sky130_fd_sc_hd__a211o_2
XFILLER_0_35_1159 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12631_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[47\] _07668_ keymem.key_mem\[6\]\[47\]
+ _07818_ _08187_ sky130_fd_sc_hd__a22o_2
X_24617_ VGND VPWR VPWR VGND clk _01110_ reset_n keymem.key_mem\[8\]\[98\] sky130_fd_sc_hd__dfrtp_2
X_21829_ VGND VPWR _01638_ _06386_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_13_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25597_ VGND VPWR VPWR VGND clk _02090_ reset_n keymem.key_mem\[0\]\[54\] sky130_fd_sc_hd__dfrtp_2
X_15350_ VPWR VGND VPWR VGND _10810_ _10811_ _10812_ _10807_ _10808_ sky130_fd_sc_hd__or4b_2
XFILLER_0_87_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12562_ VGND VPWR _08124_ _07644_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24548_ VGND VPWR VPWR VGND clk _01041_ reset_n keymem.key_mem\[8\]\[29\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14301_ VPWR VGND VPWR VGND _09770_ _09771_ _09458_ _09459_ sky130_fd_sc_hd__or3b_2
XFILLER_0_266_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15281_ VGND VPWR VGND VPWR keylen _10739_ _10740_ _10741_ _10744_ sky130_fd_sc_hd__a31o_2
XFILLER_0_48_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24479_ VGND VPWR VPWR VGND clk _00972_ reset_n keymem.key_mem\[9\]\[88\] sky130_fd_sc_hd__dfrtp_2
X_12493_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[34\] _07565_ keymem.key_mem\[4\]\[34\]
+ _07551_ _08062_ sky130_fd_sc_hd__a22o_2
XFILLER_0_123_314 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_266_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17020_ VGND VPWR VGND VPWR _03142_ _02647_ _03144_ _03143_ sky130_fd_sc_hd__a21oi_2
X_14232_ _09701_ _09703_ _09700_ _09702_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_262_1338 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_184_1196 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_21_323 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_61_492 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14163_ VGND VPWR VPWR VGND _09523_ _09634_ _09632_ _09630_ _09631_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_81_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13114_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[94\] _08577_ _08622_ _08618_ _08623_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_221_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14094_ VGND VPWR _09565_ _09354_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18971_ VPWR VGND _04805_ _04804_ enc_block.round_key\[54\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_219_930 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_197_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_195_2_Left_666 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17922_ VGND VPWR VGND VPWR _03476_ keymem.prev_key1_reg\[98\] _03879_ _03818_ sky130_fd_sc_hd__a21bo_2
X_13045_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[88\] _07872_ keymem.key_mem\[6\]\[88\]
+ _07639_ _08560_ sky130_fd_sc_hd__a22o_2
XFILLER_0_56_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdec_block block[0] block[100] block[101] block[102] block[103] block[104] block[105]
+ block[106] block[107] block[108] block[109] block[10] block[110] block[111] block[112]
+ block[113] block[114] block[115] block[116] block[117] block[118] block[119] block[11]
+ block[120] block[121] block[122] block[123] block[124] block[125] block[126] block[127]
+ block[12] block[13] block[14] block[15] block[16] block[17] block[18] block[19]
+ block[1] block[20] block[21] block[22] block[23] block[24] block[25] block[26] block[27]
+ block[28] block[29] block[2] block[30] block[31] block[32] block[33] block[34] block[35]
+ block[36] block[37] block[38] block[39] block[3] block[40] block[41] block[42] block[43]
+ block[44] block[45] block[46] block[47] block[48] block[49] block[4] block[50] block[51]
+ block[52] block[53] block[54] block[55] block[56] block[57] block[58] block[59]
+ block[5] block[60] block[61] block[62] block[63] block[64] block[65] block[66] block[67]
+ block[68] block[69] block[6] block[70] block[71] block[72] block[73] block[74] block[75]
+ block[76] block[77] block[78] block[79] block[7] block[80] block[81] block[82] block[83]
+ block[84] block[85] block[86] block[87] block[88] block[89] block[8] block[90] block[91]
+ block[92] block[93] block[94] block[95] block[96] block[97] block[98] block[99]
+ block[9] clk keylen dec_new_block\[0\] dec_new_block\[100\] dec_new_block\[101\]
+ dec_new_block\[102\] dec_new_block\[103\] dec_new_block\[104\] dec_new_block\[105\]
+ dec_new_block\[106\] dec_new_block\[107\] dec_new_block\[108\] dec_new_block\[109\]
+ dec_new_block\[10\] dec_new_block\[110\] dec_new_block\[111\] dec_new_block\[112\]
+ dec_new_block\[113\] dec_new_block\[114\] dec_new_block\[115\] dec_new_block\[116\]
+ dec_new_block\[117\] dec_new_block\[118\] dec_new_block\[119\] dec_new_block\[11\]
+ dec_new_block\[120\] dec_new_block\[121\] dec_new_block\[122\] dec_new_block\[123\]
+ dec_new_block\[124\] dec_new_block\[125\] dec_new_block\[126\] dec_new_block\[127\]
+ dec_new_block\[12\] dec_new_block\[13\] dec_new_block\[14\] dec_new_block\[15\]
+ dec_new_block\[16\] dec_new_block\[17\] dec_new_block\[18\] dec_new_block\[19\]
+ dec_new_block\[1\] dec_new_block\[20\] dec_new_block\[21\] dec_new_block\[22\] dec_new_block\[23\]
+ dec_new_block\[24\] dec_new_block\[25\] dec_new_block\[26\] dec_new_block\[27\]
+ dec_new_block\[28\] dec_new_block\[29\] dec_new_block\[2\] dec_new_block\[30\] dec_new_block\[31\]
+ dec_new_block\[32\] dec_new_block\[33\] dec_new_block\[34\] dec_new_block\[35\]
+ dec_new_block\[36\] dec_new_block\[37\] dec_new_block\[38\] dec_new_block\[39\]
+ dec_new_block\[3\] dec_new_block\[40\] dec_new_block\[41\] dec_new_block\[42\] dec_new_block\[43\]
+ dec_new_block\[44\] dec_new_block\[45\] dec_new_block\[46\] dec_new_block\[47\]
+ dec_new_block\[48\] dec_new_block\[49\] dec_new_block\[4\] dec_new_block\[50\] dec_new_block\[51\]
+ dec_new_block\[52\] dec_new_block\[53\] dec_new_block\[54\] dec_new_block\[55\]
+ dec_new_block\[56\] dec_new_block\[57\] dec_new_block\[58\] dec_new_block\[59\]
+ dec_new_block\[5\] dec_new_block\[60\] dec_new_block\[61\] dec_new_block\[62\] dec_new_block\[63\]
+ dec_new_block\[64\] dec_new_block\[65\] dec_new_block\[66\] dec_new_block\[67\]
+ dec_new_block\[68\] dec_new_block\[69\] dec_new_block\[6\] dec_new_block\[70\] dec_new_block\[71\]
+ dec_new_block\[72\] dec_new_block\[73\] dec_new_block\[74\] dec_new_block\[75\]
+ dec_new_block\[76\] dec_new_block\[77\] dec_new_block\[78\] dec_new_block\[79\]
+ dec_new_block\[7\] dec_new_block\[80\] dec_new_block\[81\] dec_new_block\[82\] dec_new_block\[83\]
+ dec_new_block\[84\] dec_new_block\[85\] dec_new_block\[86\] dec_new_block\[87\]
+ dec_new_block\[88\] dec_new_block\[89\] dec_new_block\[8\] dec_new_block\[90\] dec_new_block\[91\]
+ dec_new_block\[92\] dec_new_block\[93\] dec_new_block\[94\] dec_new_block\[95\]
+ dec_new_block\[96\] dec_new_block\[97\] dec_new_block\[98\] dec_new_block\[99\]
+ dec_new_block\[9\] dec_next dec_ready reset_n dec_round_nr\[0\] dec_round_nr\[1\]
+ dec_round_nr\[2\] dec_round_nr\[3\] enc_block.round_key\[0\] enc_block.round_key\[100\]
+ enc_block.round_key\[101\] enc_block.round_key\[102\] enc_block.round_key\[103\]
+ enc_block.round_key\[104\] enc_block.round_key\[105\] enc_block.round_key\[106\]
+ enc_block.round_key\[107\] enc_block.round_key\[108\] enc_block.round_key\[109\]
+ enc_block.round_key\[10\] enc_block.round_key\[110\] enc_block.round_key\[111\]
+ enc_block.round_key\[112\] enc_block.round_key\[113\] enc_block.round_key\[114\]
+ enc_block.round_key\[115\] enc_block.round_key\[116\] enc_block.round_key\[117\]
+ enc_block.round_key\[118\] enc_block.round_key\[119\] enc_block.round_key\[11\]
+ enc_block.round_key\[120\] enc_block.round_key\[121\] enc_block.round_key\[122\]
+ enc_block.round_key\[123\] enc_block.round_key\[124\] enc_block.round_key\[125\]
+ enc_block.round_key\[126\] enc_block.round_key\[127\] enc_block.round_key\[12\]
+ enc_block.round_key\[13\] enc_block.round_key\[14\] enc_block.round_key\[15\] enc_block.round_key\[16\]
+ enc_block.round_key\[17\] enc_block.round_key\[18\] enc_block.round_key\[19\] enc_block.round_key\[1\]
+ enc_block.round_key\[20\] enc_block.round_key\[21\] enc_block.round_key\[22\] enc_block.round_key\[23\]
+ enc_block.round_key\[24\] enc_block.round_key\[25\] enc_block.round_key\[26\] enc_block.round_key\[27\]
+ enc_block.round_key\[28\] enc_block.round_key\[29\] enc_block.round_key\[2\] enc_block.round_key\[30\]
+ enc_block.round_key\[31\] enc_block.round_key\[32\] enc_block.round_key\[33\] enc_block.round_key\[34\]
+ enc_block.round_key\[35\] enc_block.round_key\[36\] enc_block.round_key\[37\] enc_block.round_key\[38\]
+ enc_block.round_key\[39\] enc_block.round_key\[3\] enc_block.round_key\[40\] enc_block.round_key\[41\]
+ enc_block.round_key\[42\] enc_block.round_key\[43\] enc_block.round_key\[44\] enc_block.round_key\[45\]
+ enc_block.round_key\[46\] enc_block.round_key\[47\] enc_block.round_key\[48\] enc_block.round_key\[49\]
+ enc_block.round_key\[4\] enc_block.round_key\[50\] enc_block.round_key\[51\] enc_block.round_key\[52\]
+ enc_block.round_key\[53\] enc_block.round_key\[54\] enc_block.round_key\[55\] enc_block.round_key\[56\]
+ enc_block.round_key\[57\] enc_block.round_key\[58\] enc_block.round_key\[59\] enc_block.round_key\[5\]
+ enc_block.round_key\[60\] enc_block.round_key\[61\] enc_block.round_key\[62\] enc_block.round_key\[63\]
+ enc_block.round_key\[64\] enc_block.round_key\[65\] enc_block.round_key\[66\] enc_block.round_key\[67\]
+ enc_block.round_key\[68\] enc_block.round_key\[69\] enc_block.round_key\[6\] enc_block.round_key\[70\]
+ enc_block.round_key\[71\] enc_block.round_key\[72\] enc_block.round_key\[73\] enc_block.round_key\[74\]
+ enc_block.round_key\[75\] enc_block.round_key\[76\] enc_block.round_key\[77\] enc_block.round_key\[78\]
+ enc_block.round_key\[79\] enc_block.round_key\[7\] enc_block.round_key\[80\] enc_block.round_key\[81\]
+ enc_block.round_key\[82\] enc_block.round_key\[83\] enc_block.round_key\[84\] enc_block.round_key\[85\]
+ enc_block.round_key\[86\] enc_block.round_key\[87\] enc_block.round_key\[88\] enc_block.round_key\[89\]
+ enc_block.round_key\[8\] enc_block.round_key\[90\] enc_block.round_key\[91\] enc_block.round_key\[92\]
+ enc_block.round_key\[93\] enc_block.round_key\[94\] enc_block.round_key\[95\] enc_block.round_key\[96\]
+ enc_block.round_key\[97\] enc_block.round_key\[98\] enc_block.round_key\[99\] enc_block.round_key\[9\]
+ VPWR VGND aes_decipher_block
XFILLER_0_158_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17853_ VGND VPWR VPWR VGND _03814_ _03831_ keymem.prev_key0_reg\[76\] _03832_ sky130_fd_sc_hd__mux2_2
XFILLER_0_94_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16804_ VPWR VGND VGND VPWR _02947_ _10384_ _10655_ _02948_ sky130_fd_sc_hd__nor3_2
XFILLER_0_238_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14996_ VPWR VGND VGND VPWR _10459_ _10460_ _10455_ sky130_fd_sc_hd__nor2_2
X_17784_ VGND VPWR _00195_ _03784_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_88_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_234_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19523_ VPWR VGND keymem.key_mem\[12\]\[57\] _05162_ _05158_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13947_ VGND VPWR _09419_ _09418_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_233_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16735_ VGND VPWR _00045_ _02885_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_199_892 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_92_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16666_ _10243_ _02820_ keymem.round_ctr_reg\[0\] _10261_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_19454_ VPWR VGND keymem.key_mem\[12\]\[25\] _05125_ _05116_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13878_ VGND VPWR _09350_ _09349_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_134_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15617_ VGND VPWR VGND VPWR _10509_ _10594_ _10682_ _10604_ _11075_ sky130_fd_sc_hd__o22a_2
X_18405_ VPWR VGND VPWR VGND _04296_ _04054_ _04295_ sky130_fd_sc_hd__or2_2
X_12829_ VGND VPWR VGND VPWR _07691_ keymem.key_mem\[3\]\[66\] _08361_ _08363_ _08366_
+ _08365_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_29_434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19385_ VGND VPWR _00496_ _05084_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16597_ VGND VPWR VPWR VGND _11109_ _02753_ key[27] _02754_ sky130_fd_sc_hd__mux2_2
XFILLER_0_31_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1057 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_118_119 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15548_ VPWR VGND VGND VPWR _10751_ _10867_ _10569_ _10575_ _11007_ _11006_ sky130_fd_sc_hd__o221a_2
X_18336_ VGND VPWR _04234_ enc_block.block_w3_reg\[0\] _04140_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_56_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_227_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18267_ VGND VPWR _04171_ _03977_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15479_ VGND VPWR VGND VPWR _10600_ _10939_ _10937_ _10938_ _10936_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_112_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_245_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17218_ VGND VPWR VPWR VGND _03296_ keymem.key_mem\[14\]\[79\] _03322_ _03323_ sky130_fd_sc_hd__mux2_2
X_18198_ VPWR VGND VPWR VGND _04108_ _04040_ _04106_ enc_block.block_w0_reg\[11\]
+ _04097_ _00285_ sky130_fd_sc_hd__a221o_2
XFILLER_0_206_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17149_ VGND VPWR _00084_ _03260_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_13_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20160_ VGND VPWR VPWR VGND _05493_ _03492_ keymem.key_mem\[10\]\[100\] _05500_ sky130_fd_sc_hd__mux2_2
XFILLER_0_12_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_102_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20091_ VGND VPWR VPWR VGND _05457_ _03217_ keymem.key_mem\[10\]\[67\] _05464_ sky130_fd_sc_hd__mux2_2
XFILLER_0_256_579 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_239_1318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1078 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23850_ VGND VPWR VPWR VGND clk _00343_ reset_n enc_block.block_w2_reg\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_252_752 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_100_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22801_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[102\] _06858_ _06857_ _05037_ _02138_
+ sky130_fd_sc_hd__a22o_2
X_23781_ VGND VPWR VPWR VGND clk _00274_ reset_n enc_block.block_w0_reg\[0\] sky130_fd_sc_hd__dfrtp_2
X_20993_ VGND VPWR VPWR VGND _05934_ _05043_ keymem.key_mem\[7\]\[105\] _05944_ sky130_fd_sc_hd__mux2_2
XFILLER_0_174_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25520_ VGND VPWR VPWR VGND clk _02013_ reset_n keymem.key_mem\[1\]\[105\] sky130_fd_sc_hd__dfrtp_2
X_22732_ VGND VPWR VPWR VGND _06822_ keymem.key_mem\[0\]\[61\] _03162_ _06831_ sky130_fd_sc_hd__mux2_2
XFILLER_0_79_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_149_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_1468 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_250_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_149_244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_94_326 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25451_ VGND VPWR VPWR VGND clk _01944_ reset_n keymem.key_mem\[1\]\[36\] sky130_fd_sc_hd__dfrtp_2
X_22663_ VGND VPWR VPWR VGND _06798_ keymem.key_mem\[0\]\[20\] _02480_ _06803_ sky130_fd_sc_hd__mux2_2
XFILLER_0_34_1170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24402_ VGND VPWR VPWR VGND clk _00895_ reset_n keymem.key_mem\[9\]\[11\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_702 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21614_ VGND VPWR VPWR VGND _06263_ _10976_ keymem.key_mem\[4\]\[12\] _06274_ sky130_fd_sc_hd__mux2_2
X_25382_ VGND VPWR VPWR VGND clk _01875_ reset_n keymem.key_mem\[2\]\[95\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_1411 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22594_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[106\] _06775_ _06774_ _05045_ _02014_
+ sky130_fd_sc_hd__a22o_2
X_24333_ VGND VPWR VPWR VGND clk _00826_ reset_n keymem.key_mem\[10\]\[70\] sky130_fd_sc_hd__dfrtp_2
X_21545_ VGND VPWR _01504_ _06236_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_779 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_662 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_971 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_22_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24264_ VGND VPWR VPWR VGND clk _00757_ reset_n keymem.key_mem\[10\]\[1\] sky130_fd_sc_hd__dfrtp_2
X_21476_ VGND VPWR _06200_ _03287_ _01471_ _06114_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_23215_ VGND VPWR _07105_ enc_block.round_key\[1\] _07104_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20427_ VGND VPWR VPWR VGND _05638_ _03474_ keymem.key_mem\[9\]\[97\] _05642_ sky130_fd_sc_hd__mux2_2
XFILLER_0_15_194 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24195_ VGND VPWR VPWR VGND clk _00688_ reset_n keymem.key_mem\[11\]\[60\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_31_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23146_ VGND VPWR VGND VPWR _02285_ _07056_ _07010_ keymem.prev_key1_reg\[108\] sky130_fd_sc_hd__o21a_2
X_20358_ VGND VPWR VPWR VGND _05602_ _03194_ keymem.key_mem\[9\]\[64\] _05606_ sky130_fd_sc_hd__mux2_2
XFILLER_0_261_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_78_1_Right_679 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23077_ VGND VPWR VPWR VGND _07013_ keylen _07014_ _06926_ _03345_ sky130_fd_sc_hd__o211a_2
X_20289_ VGND VPWR VPWR VGND _05569_ _02862_ keymem.key_mem\[9\]\[31\] _05570_ sky130_fd_sc_hd__mux2_2
X_22028_ VGND VPWR _01728_ _06495_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_264_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_741 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14850_ VGND VPWR VGND VPWR _10296_ _10315_ _10311_ _10314_ _10306_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13801_ VGND VPWR _09273_ _08951_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14781_ VGND VPWR VGND VPWR _10247_ _10246_ _10116_ _09493_ sky130_fd_sc_hd__and3b_2
X_23979_ VGND VPWR VPWR VGND clk _00472_ reset_n keymem.key_mem\[13\]\[100\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_202_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11993_ VGND VPWR _07596_ _07595_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_192_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16520_ VPWR VGND VPWR VGND _02680_ keymem.prev_key1_reg\[88\] sky130_fd_sc_hd__inv_2
X_13732_ VGND VPWR _09204_ _09203_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25718_ keymem.prev_key1_reg\[34\] clk _02211_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_58_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_97_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16451_ VGND VPWR VGND VPWR _11610_ _02611_ _02612_ _11481_ _02417_ sky130_fd_sc_hd__nor4_2
X_13663_ VPWR VGND VPWR VGND _09044_ _09005_ _08991_ _08977_ _09135_ sky130_fd_sc_hd__or4_2
X_25649_ VGND VPWR VPWR VGND clk _02142_ reset_n keymem.key_mem\[0\]\[106\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_210_170 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15402_ VPWR VGND VGND VPWR _10588_ _10863_ _10633_ sky130_fd_sc_hd__nor2_2
X_19170_ VGND VPWR VPWR VGND _04928_ _04947_ keymem.key_mem\[13\]\[46\] _04948_ sky130_fd_sc_hd__mux2_2
X_12614_ VGND VPWR VGND VPWR _08172_ _07839_ keymem.key_mem\[11\]\[45\] _08169_ _08171_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_155_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16382_ VGND VPWR VGND VPWR _02543_ _02542_ _02545_ _02544_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_213_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13594_ VPWR VGND VPWR VGND _09031_ _09065_ _08971_ _09009_ _09066_ sky130_fd_sc_hd__or4_2
XFILLER_0_26_415 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_53_201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18121_ VPWR VGND VPWR VGND _04037_ block[101] _03980_ enc_block.block_w3_reg\[5\]
+ _04007_ _04038_ sky130_fd_sc_hd__a221o_2
XFILLER_0_186_1236 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15333_ VPWR VGND VPWR VGND _10689_ _10794_ _10795_ _10605_ _10622_ sky130_fd_sc_hd__or4b_2
XFILLER_0_108_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12545_ VGND VPWR VGND VPWR _08016_ keymem.key_mem\[7\]\[39\] _08106_ _08108_ _08109_
+ _08069_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_48_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18052_ VGND VPWR _03974_ _03973_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15264_ VPWR VGND VPWR VGND _10631_ _10726_ _10724_ _10471_ _10727_ sky130_fd_sc_hd__or4_2
XFILLER_0_227_1233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12476_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[33\] _07902_ keymem.key_mem\[10\]\[33\]
+ _07785_ _08046_ sky130_fd_sc_hd__a22o_2
X_17003_ VGND VPWR VGND VPWR _03129_ _11151_ key[186] _03123_ _03128_ sky130_fd_sc_hd__a211o_2
X_14215_ VGND VPWR VGND VPWR _09686_ _09685_ _09682_ _09681_ _09680_ sky130_fd_sc_hd__and4_2
XFILLER_0_46_1030 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15195_ VGND VPWR VGND VPWR _10190_ _10189_ _10658_ _10655_ _10659_ sky130_fd_sc_hd__a31o_2
XFILLER_0_240_1411 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14146_ VPWR VGND VGND VPWR _09434_ _09617_ _09335_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_256_Right_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18954_ VPWR VGND VPWR VGND _04789_ _04788_ _04787_ enc_block.block_w2_reg\[20\]
+ _04709_ _00360_ sky130_fd_sc_hd__a221o_2
X_14077_ VGND VPWR VGND VPWR _09545_ _08927_ _09548_ _09547_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_67_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13028_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[86\] _07760_ keymem.key_mem\[9\]\[86\]
+ _07672_ _08545_ sky130_fd_sc_hd__a22o_2
X_17905_ VGND VPWR VGND VPWR _03730_ keymem.prev_key0_reg\[92\] _03867_ _03432_ _00233_
+ sky130_fd_sc_hd__a2bb2o_2
X_18885_ VGND VPWR _04727_ enc_block.block_w0_reg\[13\] _04656_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17836_ VGND VPWR _00211_ _03820_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_177_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_59_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_774 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_571 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_234_1226 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_233_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17767_ VGND VPWR _00188_ _03774_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14979_ VGND VPWR _10443_ _10442_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_171_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19506_ VGND VPWR VPWR VGND _05151_ _04953_ keymem.key_mem\[12\]\[49\] _05153_ sky130_fd_sc_hd__mux2_2
XFILLER_0_178_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16718_ VGND VPWR VGND VPWR _09530_ _09529_ _02870_ _02869_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_88_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17698_ VGND VPWR _03729_ _03728_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_53_1056 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19437_ VGND VPWR VGND VPWR _05115_ keymem.key_mem_we _11547_ _05109_ _00517_ sky130_fd_sc_hd__a31o_2
X_16649_ VGND VPWR VGND VPWR _02802_ keymem.prev_key1_reg\[93\] _02804_ _02801_ sky130_fd_sc_hd__nand3_2
XFILLER_0_14_1029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_123_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_169_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19368_ VPWR VGND keymem.key_mem_we _05073_ _03613_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_18_938 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18319_ VGND VPWR VGND VPWR _04217_ _04216_ _04219_ _04215_ sky130_fd_sc_hd__a21oi_2
X_19299_ VGND VPWR _00468_ _05026_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_114_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21330_ VGND VPWR VPWR VGND _06117_ _10283_ keymem.key_mem\[5\]\[6\] _06124_ sky130_fd_sc_hd__mux2_2
XFILLER_0_5_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21261_ VGND VPWR VPWR VGND _06076_ _03511_ keymem.key_mem\[6\]\[103\] _06086_ sky130_fd_sc_hd__mux2_2
X_23000_ VGND VPWR _02228_ _06967_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20212_ VGND VPWR VPWR VGND _05388_ _03654_ keymem.key_mem\[10\]\[125\] _05527_ sky130_fd_sc_hd__mux2_2
XFILLER_0_40_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21192_ VGND VPWR VPWR VGND _06040_ _03245_ keymem.key_mem\[6\]\[70\] _06050_ sky130_fd_sc_hd__mux2_2
XFILLER_0_106_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20143_ VGND VPWR VPWR VGND _05482_ _03435_ keymem.key_mem\[10\]\[92\] _05491_ sky130_fd_sc_hd__mux2_2
XFILLER_0_25_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20074_ VGND VPWR VPWR VGND _05446_ _03140_ keymem.key_mem\[10\]\[59\] _05455_ sky130_fd_sc_hd__mux2_2
X_24951_ VGND VPWR VPWR VGND clk _01444_ reset_n keymem.key_mem\[5\]\[48\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_244_549 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23902_ VGND VPWR VPWR VGND clk _00395_ reset_n keymem.key_mem\[13\]\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24882_ VGND VPWR VPWR VGND clk _01375_ reset_n keymem.key_mem\[6\]\[107\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_225_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23833_ VGND VPWR VPWR VGND clk _00326_ reset_n enc_block.block_w1_reg\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_252_582 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_217_1446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_169_317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_217_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23764_ keymem.prev_key0_reg\[120\] clk _00261_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20976_ VGND VPWR _01236_ _05935_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25503_ VGND VPWR VPWR VGND clk _01996_ reset_n keymem.key_mem\[1\]\[88\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_67_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22715_ VGND VPWR _02087_ _06823_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_177_361 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_67_359 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23695_ keymem.prev_key0_reg\[51\] clk _00192_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_14_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25434_ VGND VPWR VPWR VGND clk _01927_ reset_n keymem.key_mem\[1\]\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_36_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22646_ VGND VPWR VPWR VGND _06785_ keymem.key_mem\[0\]\[12\] _10977_ _06794_ sky130_fd_sc_hd__mux2_2
XFILLER_0_63_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25365_ VGND VPWR VPWR VGND clk _01858_ reset_n keymem.key_mem\[2\]\[78\] sky130_fd_sc_hd__dfrtp_2
X_22577_ VGND VPWR VPWR VGND _06701_ keymem.key_mem\[1\]\[93\] _03444_ _06772_ sky130_fd_sc_hd__mux2_2
XFILLER_0_183_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_114_1_Left_381 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24316_ VGND VPWR VPWR VGND clk _00809_ reset_n keymem.key_mem\[10\]\[53\] sky130_fd_sc_hd__dfrtp_2
X_12330_ VGND VPWR _07913_ _07550_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21528_ VGND VPWR _01496_ _06227_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_228_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25296_ VGND VPWR VPWR VGND clk _01789_ reset_n keymem.key_mem\[2\]\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_259_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12261_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[15\] _07703_ keymem.key_mem\[14\]\[15\]
+ _07782_ _07849_ sky130_fd_sc_hd__a22o_2
X_24247_ VGND VPWR VPWR VGND clk _00740_ reset_n keymem.key_mem\[11\]\[112\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_105_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21459_ VGND VPWR _01463_ _06191_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_146_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14000_ VPWR VGND VGND VPWR _09247_ _09472_ _09361_ sky130_fd_sc_hd__nor2_2
XFILLER_0_32_974 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_1214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12192_ VGND VPWR _07785_ _07742_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24178_ VGND VPWR VPWR VGND clk _00671_ reset_n keymem.key_mem\[11\]\[43\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_31_495 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23129_ VPWR VGND VPWR VGND _07045_ keymem.prev_key1_reg\[103\] _06878_ sky130_fd_sc_hd__or2_2
XFILLER_0_43_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_372 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_247_387 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15951_ VGND VPWR VGND VPWR _11407_ _11229_ _11228_ _11272_ _11288_ sky130_fd_sc_hd__and4_2
XFILLER_0_37_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14902_ VGND VPWR VGND VPWR _10367_ _10366_ _10364_ _10363_ _10330_ sky130_fd_sc_hd__o211ai_2
X_15882_ VGND VPWR _11338_ _11258_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18670_ VPWR VGND _04534_ _04533_ enc_block.round_key\[88\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_250_519 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_235_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_204_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17621_ VGND VPWR VPWR VGND _03675_ _03671_ keymem.prev_key0_reg\[0\] _03676_ sky130_fd_sc_hd__mux2_2
X_14833_ VGND VPWR VGND VPWR _09480_ _09475_ _09349_ _09450_ _10298_ sky130_fd_sc_hd__o22a_2
XFILLER_0_192_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_958 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_144_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14764_ _10215_ _10230_ keymem.round_ctr_reg\[0\] _10229_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_17552_ VGND VPWR VGND VPWR _03616_ _10328_ _02877_ key[120] sky130_fd_sc_hd__o21a_2
X_11976_ VGND VPWR _07579_ _07578_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_114_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_224_40 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_187_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13715_ VGND VPWR VGND VPWR _09186_ _09153_ _09187_ _09056_ sky130_fd_sc_hd__a21oi_2
X_16503_ VGND VPWR _00035_ _02663_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_233_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17483_ VGND VPWR _00122_ _03556_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_168_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14695_ VPWR VGND VPWR VGND _10160_ _10161_ _10162_ _09801_ _10157_ sky130_fd_sc_hd__or4b_2
XFILLER_0_230_298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_1141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19222_ VGND VPWR _04979_ _04879_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_2_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13646_ VPWR VGND VPWR VGND _09118_ _09106_ _09107_ _09108_ _09111_ _09117_ sky130_fd_sc_hd__o311a_2
X_16434_ VGND VPWR VGND VPWR key[22] _09930_ _02595_ _02594_ _02596_ sky130_fd_sc_hd__o22a_2
XFILLER_0_6_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_510 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_629 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16365_ VGND VPWR VGND VPWR _11250_ _11298_ _02528_ _11318_ sky130_fd_sc_hd__a21oi_2
X_19153_ VGND VPWR _00412_ _04936_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13577_ VPWR VGND VPWR VGND _09013_ _09005_ _08990_ _09001_ _09049_ sky130_fd_sc_hd__or4_2
XFILLER_0_14_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15316_ VPWR VGND VGND VPWR _10488_ _10545_ _10778_ _10503_ _10635_ sky130_fd_sc_hd__o22ai_2
X_18104_ VPWR VGND _04022_ enc_block.block_w3_reg\[7\] enc_block.block_w3_reg\[3\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_12528_ VGND VPWR VGND VPWR _08094_ _08008_ keymem.key_mem\[2\]\[37\] _08091_ _08093_
+ sky130_fd_sc_hd__a211o_2
X_16296_ VGND VPWR VGND VPWR _02459_ _02412_ keymem.prev_key0_reg\[116\] _02460_ sky130_fd_sc_hd__a21o_2
XFILLER_0_136_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19084_ VGND VPWR _04896_ _04877_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_23_930 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15247_ VPWR VGND VGND VPWR _10545_ _10710_ _10526_ sky130_fd_sc_hd__nor2_2
X_18035_ VGND VPWR _03957_ _03956_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12459_ VGND VPWR VGND VPWR _07778_ keymem.key_mem\[3\]\[31\] _08028_ _08030_ _08031_
+ _07573_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_22_440 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15178_ VGND VPWR VGND VPWR _10528_ _10522_ _10642_ _10629_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_125_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_160_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_367 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14129_ VGND VPWR VGND VPWR _09333_ _09375_ _09559_ _09419_ _09600_ sky130_fd_sc_hd__o22a_2
XFILLER_0_1_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_249_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19986_ VGND VPWR VPWR VGND _05400_ _11547_ keymem.key_mem\[10\]\[17\] _05409_ sky130_fd_sc_hd__mux2_2
XFILLER_0_238_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_238_387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18937_ VGND VPWR _04774_ _04771_ _04773_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_185_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_118_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_241_508 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18868_ VGND VPWR _04712_ _04638_ _04711_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_241_519 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_158_2_Left_629 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_94_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17819_ VGND VPWR VPWR VGND _03719_ key[194] keymem.prev_key1_reg\[66\] _03808_ sky130_fd_sc_hd__mux2_2
XFILLER_0_175_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18799_ VPWR VGND VGND VPWR _04650_ _04646_ _04648_ sky130_fd_sc_hd__nand2_2
XFILLER_0_171_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20830_ VPWR VGND keymem.key_mem\[7\]\[28\] _05858_ _05856_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_49_326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_132_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20761_ VGND VPWR _01139_ _05817_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_159_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_58_860 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_119_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22500_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[49\] _06737_ _06736_ _04953_ _01957_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_18_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23480_ VGND VPWR _07342_ _04274_ _02333_ _07115_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_20692_ VGND VPWR _01106_ _05781_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22431_ VGND VPWR _01917_ _06709_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_18_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25150_ VGND VPWR VPWR VGND clk _01643_ reset_n keymem.key_mem\[4\]\[119\] sky130_fd_sc_hd__dfrtp_2
X_22362_ VGND VPWR VPWR VGND _06669_ _03533_ keymem.key_mem\[2\]\[106\] _06672_ sky130_fd_sc_hd__mux2_2
XFILLER_0_33_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24101_ VGND VPWR VPWR VGND clk _00594_ reset_n keymem.key_mem\[12\]\[94\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_182_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21313_ VPWR VGND VPWR VGND _05530_ keymem.round_ctr_reg\[2\] _06113_ keymem.round_ctr_reg\[1\]
+ keymem.round_ctr_reg\[3\] sky130_fd_sc_hd__or4b_2
XFILLER_0_245_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25081_ VGND VPWR VPWR VGND clk _01574_ reset_n keymem.key_mem\[4\]\[50\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_206_1114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_66_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22293_ VGND VPWR VPWR VGND _06634_ _03267_ keymem.key_mem\[2\]\[73\] _06636_ sky130_fd_sc_hd__mux2_2
XFILLER_0_143_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_182_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24032_ VGND VPWR VPWR VGND clk _00525_ reset_n keymem.key_mem\[12\]\[25\] sky130_fd_sc_hd__dfrtp_2
X_21244_ VGND VPWR _01362_ _06077_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_83_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_143_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_495 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_40_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21175_ VGND VPWR _01329_ _06041_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_257_663 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_245_825 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_102_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20126_ VGND VPWR _05482_ _05387_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20057_ VGND VPWR _05446_ _05388_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24934_ VGND VPWR VPWR VGND clk _01427_ reset_n keymem.key_mem\[5\]\[31\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_244_368 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_245_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_175_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24865_ VGND VPWR VPWR VGND clk _01358_ reset_n keymem.key_mem\[6\]\[90\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_193_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11830_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[18\] dec_new_block\[82\]
+ _07479_ sky130_fd_sc_hd__mux2_2
X_23816_ VGND VPWR VPWR VGND clk _00309_ reset_n enc_block.block_w1_reg\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_252_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_154_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24796_ VGND VPWR VPWR VGND clk _01289_ reset_n keymem.key_mem\[6\]\[21\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_90_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11761_ VGND VPWR result[47] _07444_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_261_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23747_ keymem.prev_key0_reg\[103\] clk _00244_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_67_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20959_ VGND VPWR _01228_ _05926_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_36_1084 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_51_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13500_ VGND VPWR VPWR VGND _08963_ _08971_ _08958_ _08972_ sky130_fd_sc_hd__or3_2
X_14480_ VGND VPWR VGND VPWR _09106_ _09797_ _09948_ _09828_ _09949_ sky130_fd_sc_hd__o22a_2
XFILLER_0_230_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_329 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23678_ keymem.prev_key0_reg\[34\] clk _00175_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_11692_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[13\] dec_new_block\[13\]
+ _07410_ sky130_fd_sc_hd__mux2_2
XFILLER_0_64_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13431_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[126\] _07651_ keymem.key_mem\[1\]\[126\]
+ _07670_ _08908_ sky130_fd_sc_hd__a22o_2
XFILLER_0_192_150 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25417_ VGND VPWR VPWR VGND clk _01910_ reset_n keymem.key_mem\[1\]\[2\] sky130_fd_sc_hd__dfrtp_2
X_22629_ VGND VPWR _06785_ _06784_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_3_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16150_ VGND VPWR VPWR VGND _11289_ _11273_ _11226_ _11604_ sky130_fd_sc_hd__or3_2
X_25348_ VGND VPWR VPWR VGND clk _01841_ reset_n keymem.key_mem\[2\]\[61\] sky130_fd_sc_hd__dfrtp_2
X_13362_ VPWR VGND VPWR VGND _08845_ keymem.key_mem\[8\]\[119\] _07541_ keymem.key_mem\[1\]\[119\]
+ _07671_ _08846_ sky130_fd_sc_hd__a221o_2
XFILLER_0_90_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15101_ VGND VPWR _10565_ _10449_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12313_ VGND VPWR VGND VPWR _07897_ _07877_ keymem.key_mem\[10\]\[19\] _07895_ _07896_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_180_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16081_ VGND VPWR VPWR VGND _11458_ _11533_ _11534_ _11536_ sky130_fd_sc_hd__or3_2
X_25279_ VGND VPWR VPWR VGND clk _01772_ reset_n keymem.key_mem\[3\]\[120\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_210_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13293_ VGND VPWR VGND VPWR _08784_ _07839_ keymem.key_mem\[11\]\[112\] _08781_ _08783_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_161_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15032_ VGND VPWR _10496_ _10495_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12244_ VPWR VGND VPWR VGND _07832_ keymem.key_mem\[10\]\[14\] _07629_ keymem.key_mem\[12\]\[14\]
+ _07579_ _07833_ sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_15_Left_283 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_267_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_241_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19840_ VGND VPWR _00705_ _05330_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_236_803 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12175_ VGND VPWR VGND VPWR _07547_ keymem.key_mem\[2\]\[9\] _07766_ _07768_ _07769_
+ _07616_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_248_685 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19771_ VGND VPWR _00672_ _05294_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16983_ VGND VPWR _00068_ _03110_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_262_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18722_ _04578_ _04580_ _04560_ _04579_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_257_1045 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15934_ VGND VPWR VGND VPWR _11390_ _11229_ _11289_ _11227_ _11226_ sky130_fd_sc_hd__and4_2
XFILLER_0_64_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_262_176 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18653_ VPWR VGND VPWR VGND _04518_ block[86] _04487_ enc_block.block_w2_reg\[22\]
+ _04425_ _04519_ sky130_fd_sc_hd__a221o_2
X_15865_ VGND VPWR VGND VPWR _11316_ _11284_ _11320_ _11318_ _11321_ sky130_fd_sc_hd__o22a_2
X_17604_ VGND VPWR VPWR VGND _09863_ keymem.key_mem\[14\]\[126\] _03661_ _03662_ sky130_fd_sc_hd__mux2_2
X_14816_ VGND VPWR VPWR VGND _10277_ _10272_ _10282_ _10281_ _10280_ sky130_fd_sc_hd__o211a_2
X_18584_ VPWR VGND VPWR VGND _04456_ block[79] _04330_ enc_block.block_w3_reg\[15\]
+ _04425_ _04457_ sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_24_Left_292 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15796_ VGND VPWR _11252_ _11251_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_59_635 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17535_ VGND VPWR _00129_ _03601_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_15_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14747_ VPWR VGND VGND VPWR _09132_ _09069_ _09107_ _09221_ _10213_ _10212_ sky130_fd_sc_hd__o221a_2
X_11959_ VGND VPWR _07562_ _07561_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_168_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_15_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14678_ VGND VPWR VPWR VGND _10144_ _10103_ _10102_ _10145_ sky130_fd_sc_hd__mux2_2
X_17466_ VGND VPWR VGND VPWR _03541_ _02995_ _03542_ keylen sky130_fd_sc_hd__a21oi_2
XFILLER_0_55_830 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19205_ VGND VPWR VGND VPWR _04969_ keymem.key_mem_we _03140_ _04968_ _00431_ sky130_fd_sc_hd__a31o_2
X_16417_ VPWR VGND VPWR VGND _11569_ _02432_ _11592_ _11498_ _02579_ sky130_fd_sc_hd__or4_2
X_13629_ VPWR VGND VPWR VGND _09044_ _09005_ _09045_ _09043_ _09101_ sky130_fd_sc_hd__or4_2
XFILLER_0_89_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17397_ VGND VPWR VGND VPWR _03482_ _03302_ _08937_ key[99] sky130_fd_sc_hd__o21a_2
XFILLER_0_54_351 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19136_ VGND VPWR VGND VPWR _04925_ keymem.key_mem_we _02894_ _04924_ _00406_ sky130_fd_sc_hd__a31o_2
X_16348_ VGND VPWR VGND VPWR _11316_ _11327_ _11332_ _11399_ _02511_ sky130_fd_sc_hd__o22a_2
XFILLER_0_171_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_192 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16279_ VGND VPWR VGND VPWR _11276_ _11286_ _02439_ _02440_ _02443_ _02442_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_42_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19067_ VPWR VGND keymem.key_mem\[13\]\[5\] _04886_ _04880_ VPWR VGND sky130_fd_sc_hd__and2_2
X_18018_ VGND VPWR VGND VPWR _00270_ _03943_ _03941_ enc_block.round\[1\] sky130_fd_sc_hd__o21a_2
XFILLER_0_125_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_65_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_196_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_96_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19969_ VGND VPWR _00765_ _05399_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22980_ VGND VPWR VGND VPWR _02220_ _06955_ _06954_ keymem.prev_key1_reg\[43\] sky130_fd_sc_hd__o21a_2
X_21931_ VGND VPWR VGND VPWR _06443_ keymem.key_mem_we _02862_ _06432_ _01683_ sky130_fd_sc_hd__a31o_2
XFILLER_0_218_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1095 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24650_ VGND VPWR VPWR VGND clk _01143_ reset_n keymem.key_mem\[7\]\[3\] sky130_fd_sc_hd__dfrtp_2
X_21862_ VGND VPWR _06406_ _06405_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_145_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_136_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23601_ VGND VPWR VPWR VGND clk _00102_ reset_n keymem.key_mem\[14\]\[90\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_210_736 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_72_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20813_ VGND VPWR VGND VPWR _05848_ keymem.key_mem_we _02480_ _05838_ _01160_ sky130_fd_sc_hd__a31o_2
XFILLER_0_166_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24581_ VGND VPWR VPWR VGND clk _01074_ reset_n keymem.key_mem\[8\]\[62\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21793_ VGND VPWR VPWR VGND _06366_ _03474_ keymem.key_mem\[4\]\[97\] _06368_ sky130_fd_sc_hd__mux2_2
XFILLER_0_37_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23532_ VGND VPWR VPWR VGND clk _00033_ reset_n keymem.key_mem\[14\]\[21\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20744_ VGND VPWR VPWR VGND _05805_ _03613_ keymem.key_mem\[8\]\[119\] _05809_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_114_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_107_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1509 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_275 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23463_ VPWR VGND _07327_ enc_block.block_w0_reg\[18\] enc_block.block_w2_reg\[3\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_20675_ VGND VPWR VPWR VGND _05772_ _03383_ keymem.key_mem\[8\]\[86\] _05773_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_565 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_46_874 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25202_ VGND VPWR VPWR VGND clk _01695_ reset_n keymem.key_mem\[3\]\[43\] sky130_fd_sc_hd__dfrtp_2
X_22414_ VGND VPWR _01910_ _06699_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23394_ VPWR VGND _07266_ enc_block.block_w0_reg\[18\] enc_block.block_w3_reg\[27\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_60_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25133_ VGND VPWR VPWR VGND clk _01626_ reset_n keymem.key_mem\[4\]\[102\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22345_ VGND VPWR VPWR VGND _06658_ _03480_ keymem.key_mem\[2\]\[98\] _06663_ sky130_fd_sc_hd__mux2_2
XFILLER_0_249_405 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_60_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25064_ VGND VPWR VPWR VGND clk _01557_ reset_n keymem.key_mem\[4\]\[33\] sky130_fd_sc_hd__dfrtp_2
X_22276_ VGND VPWR VPWR VGND _06622_ _03202_ keymem.key_mem\[2\]\[65\] _06627_ sky130_fd_sc_hd__mux2_2
XFILLER_0_13_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_83_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24015_ VGND VPWR VPWR VGND clk _00508_ reset_n keymem.key_mem\[12\]\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_143_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21227_ VGND VPWR _01354_ _06068_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_44_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21158_ VGND VPWR _01321_ _06032_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_218_847 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20109_ VGND VPWR _05473_ _03287_ _00831_ _05402_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_13980_ VGND VPWR VGND VPWR _09452_ _09317_ _09315_ _09319_ _09331_ sky130_fd_sc_hd__a211o_2
XFILLER_0_219_1316 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_205_508 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21089_ VGND VPWR _05996_ _05971_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12931_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[76\] _08449_ _08457_ _08453_ _08458_
+ sky130_fd_sc_hd__o22a_2
X_24917_ VGND VPWR VPWR VGND clk _01410_ reset_n keymem.key_mem\[5\]\[14\] sky130_fd_sc_hd__dfrtp_2
X_12862_ VGND VPWR enc_block.round_key\[69\] _08395_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15650_ VGND VPWR VGND VPWR _11107_ _11106_ _11105_ keymem.prev_key1_reg\[79\] _10286_
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_34_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24848_ VGND VPWR VPWR VGND clk _01341_ reset_n keymem.key_mem\[6\]\[73\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_154_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14601_ VPWR VGND VPWR VGND _10066_ _10068_ _10067_ _09880_ _10069_ sky130_fd_sc_hd__or4_2
X_11813_ VGND VPWR result[73] _07470_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_90_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15581_ VGND VPWR _11040_ _11039_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_150_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12793_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[63\] _07963_ keymem.key_mem\[4\]\[63\]
+ _07693_ _08333_ sky130_fd_sc_hd__a22o_2
XFILLER_0_205_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24779_ VGND VPWR VPWR VGND clk _01272_ reset_n keymem.key_mem\[6\]\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_55_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14532_ VPWR VGND VGND VPWR _09087_ _09108_ _10000_ _09153_ _09211_ _08999_ sky130_fd_sc_hd__o32ai_2
XFILLER_0_95_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17320_ VGND VPWR _03414_ keymem.prev_key0_reg\[90\] _02728_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_90_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11744_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[7\] dec_new_block\[39\]
+ _07436_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_279 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_189_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14463_ VGND VPWR _09932_ _09516_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17251_ VPWR VGND VGND VPWR _03352_ key[211] _10092_ sky130_fd_sc_hd__nand2_2
X_11675_ VGND VPWR result[4] _07401_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_3_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16202_ VGND VPWR VGND VPWR _11420_ _11466_ _02367_ _11469_ sky130_fd_sc_hd__a21oi_2
X_13414_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[124\] _08027_ _08892_ _08886_ _08893_
+ sky130_fd_sc_hd__o22a_2
X_17182_ VGND VPWR _03289_ _02708_ _03290_ _10969_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_14394_ VGND VPWR _09864_ _09863_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_265_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16133_ VGND VPWR VPWR VGND _11345_ _11283_ _11587_ _11586_ _11585_ sky130_fd_sc_hd__o211a_2
X_13345_ VGND VPWR enc_block.round_key\[117\] _08830_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_153_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_59_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_24_579 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_267_202 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16064_ VPWR VGND VGND VPWR _11519_ _11517_ _11518_ sky130_fd_sc_hd__nand2_2
XFILLER_0_126_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_161_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13276_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[110\] _07536_ _08768_ _08764_ enc_block.round_key\[110\]
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_122_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15015_ VPWR VGND VGND VPWR _10474_ _10462_ _10479_ _10476_ _10478_ _10475_ sky130_fd_sc_hd__o32ai_2
XFILLER_0_20_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_275 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_126_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12227_ VGND VPWR _07818_ _07759_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_161_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19823_ VGND VPWR _00697_ _05321_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12158_ VGND VPWR _07753_ _07752_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_97_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_235_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19754_ VGND VPWR _00664_ _05285_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16966_ VPWR VGND VPWR VGND _03095_ keymem.prev_key1_reg\[55\] sky130_fd_sc_hd__inv_2
X_12089_ VGND VPWR VGND VPWR _07688_ _07683_ keymem.key_mem\[5\]\[4\] _07684_ _07687_
+ sky130_fd_sc_hd__a211o_2
X_18705_ _04563_ _04565_ _04560_ _04564_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_237_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15917_ VGND VPWR VGND VPWR _11372_ _11370_ _11278_ _11257_ _11286_ _11373_ sky130_fd_sc_hd__o32a_2
XPHY_EDGE_ROW_32_Left_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19685_ VGND VPWR _00631_ _05249_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16897_ VGND VPWR VGND VPWR _11155_ _11154_ _03033_ _03032_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_56_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18636_ VPWR VGND VPWR VGND _04503_ _04459_ _04502_ enc_block.block_w1_reg\[20\]
+ _04424_ _00328_ sky130_fd_sc_hd__a221o_2
XFILLER_0_257_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15848_ VPWR VGND VPWR VGND _11264_ _11216_ _11243_ _11232_ _11304_ sky130_fd_sc_hd__or4_2
XFILLER_0_133_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18567_ VGND VPWR VPWR VGND _04316_ enc_block.block_w1_reg\[13\] _04125_ _04442_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_73_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15779_ VGND VPWR _11235_ _11234_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_34_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_169_1_Right_770 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_148_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_231_1059 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17518_ VGND VPWR _00127_ _03586_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_34_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18498_ VGND VPWR _04380_ _04314_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_213_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17449_ VGND VPWR _03527_ _09543_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_131_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_15_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20460_ VGND VPWR VPWR VGND _05649_ _03573_ keymem.key_mem\[9\]\[113\] _05659_ sky130_fd_sc_hd__mux2_2
XFILLER_0_171_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_54_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19119_ VGND VPWR _04915_ _04879_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_6_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20391_ VGND VPWR VPWR VGND _05614_ _03330_ keymem.key_mem\[9\]\[80\] _05623_ sky130_fd_sc_hd__mux2_2
XFILLER_0_42_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22130_ VGND VPWR _01777_ _06548_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_144_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Right_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_112_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_590 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_80_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_140_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1050 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22061_ VGND VPWR VGND VPWR _06512_ keymem.key_mem_we _03435_ _06498_ _01744_ sky130_fd_sc_hd__a31o_2
XFILLER_0_80_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_11_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21012_ VGND VPWR VPWR VGND _05945_ _05062_ keymem.key_mem\[7\]\[114\] _05954_ sky130_fd_sc_hd__mux2_2
XFILLER_0_220_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_215_806 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25820_ VGND VPWR VPWR VGND clk _02313_ reset_n enc_block.block_w3_reg\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_255_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_220_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25751_ keymem.prev_key1_reg\[67\] clk _02244_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_255_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22963_ VGND VPWR VGND VPWR _06888_ _06944_ _02213_ _06945_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_123_1_Left_390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24702_ VGND VPWR VPWR VGND clk _01195_ reset_n keymem.key_mem\[7\]\[55\] sky130_fd_sc_hd__dfrtp_2
X_21914_ VGND VPWR VGND VPWR _06434_ keymem.key_mem_we _02661_ _06432_ _01675_ sky130_fd_sc_hd__a31o_2
X_25682_ VGND VPWR VPWR VGND clk _02175_ reset_n keymem.round_ctr_reg\[3\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_21_Right_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22894_ VGND VPWR _02187_ _06902_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_151_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1284 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_214_1235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24633_ VGND VPWR VPWR VGND clk _01126_ reset_n keymem.key_mem\[8\]\[114\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_139_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21845_ VGND VPWR VPWR VGND _06388_ _03633_ keymem.key_mem\[4\]\[122\] _06395_ sky130_fd_sc_hd__mux2_2
XFILLER_0_151_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24564_ VGND VPWR VPWR VGND clk _01057_ reset_n keymem.key_mem\[8\]\[45\] sky130_fd_sc_hd__dfrtp_2
X_21776_ VGND VPWR VPWR VGND _06355_ _03409_ keymem.key_mem\[4\]\[89\] _06359_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23515_ VGND VPWR VPWR VGND clk _00016_ reset_n keymem.key_mem\[14\]\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20727_ VGND VPWR VPWR VGND _05794_ _03560_ keymem.key_mem\[8\]\[111\] _05800_ sky130_fd_sc_hd__mux2_2
X_24495_ VGND VPWR VPWR VGND clk _00988_ reset_n keymem.key_mem\[9\]\[104\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_276 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_135_345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_142_1_Left_409 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23446_ VGND VPWR _07312_ enc_block.block_w0_reg\[17\] _07097_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20658_ VGND VPWR VPWR VGND _05761_ _03314_ keymem.key_mem\[8\]\[78\] _05764_ sky130_fd_sc_hd__mux2_2
XFILLER_0_262_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23377_ VPWR VGND VPWR VGND _07251_ _07247_ _07249_ sky130_fd_sc_hd__or2_2
XFILLER_0_21_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20589_ VGND VPWR VPWR VGND _05725_ _03006_ keymem.key_mem\[8\]\[45\] _05728_ sky130_fd_sc_hd__mux2_2
XFILLER_0_225_1320 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25116_ VGND VPWR VPWR VGND clk _01609_ reset_n keymem.key_mem\[4\]\[85\] sky130_fd_sc_hd__dfrtp_2
X_13130_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[96\] _07579_ keymem.key_mem\[8\]\[96\]
+ _07753_ _08637_ sky130_fd_sc_hd__a22o_2
X_22328_ VGND VPWR VPWR VGND _06647_ _03417_ keymem.key_mem\[2\]\[90\] _06654_ sky130_fd_sc_hd__mux2_2
XFILLER_0_267_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13061_ VGND VPWR VGND VPWR _08575_ _07731_ keymem.key_mem\[13\]\[89\] _08572_ _08574_
+ sky130_fd_sc_hd__a211o_2
X_25047_ VGND VPWR VPWR VGND clk _01540_ reset_n keymem.key_mem\[4\]\[16\] sky130_fd_sc_hd__dfrtp_2
X_22259_ VGND VPWR VPWR VGND _06611_ _03118_ keymem.key_mem\[2\]\[57\] _06618_ sky130_fd_sc_hd__mux2_2
XFILLER_0_108_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12012_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[1\] _07564_ keymem.key_mem\[8\]\[1\]
+ _07539_ _07614_ sky130_fd_sc_hd__a22o_2
XFILLER_0_79_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_452 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16820_ VGND VPWR VGND VPWR keylen _02963_ _02962_ keymem.prev_key1_reg\[41\] _10739_
+ _10740_ sky130_fd_sc_hd__a311oi_2
X_16751_ VGND VPWR VGND VPWR _02900_ _09721_ _09719_ key[35] sky130_fd_sc_hd__o21a_2
XFILLER_0_232_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13963_ VGND VPWR VGND VPWR _09431_ _09425_ _09398_ _09434_ _09435_ sky130_fd_sc_hd__a31o_2
XFILLER_0_45_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15702_ VGND VPWR VGND VPWR _11155_ _11154_ _11158_ _11157_ sky130_fd_sc_hd__a21oi_2
X_19470_ VGND VPWR _00532_ _05133_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12914_ VPWR VGND VPWR VGND _08441_ keymem.key_mem\[5\]\[75\] _07811_ keymem.key_mem\[9\]\[75\]
+ _07738_ _08442_ sky130_fd_sc_hd__a221o_2
X_13894_ VGND VPWR _09366_ _09365_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16682_ VPWR VGND VPWR VGND _02836_ key[158] _10286_ sky130_fd_sc_hd__or2_2
X_18421_ VGND VPWR _04309_ _04306_ _04308_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15633_ VGND VPWR _11090_ keymem.round_ctr_reg\[0\] _11091_ _11057_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_119_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12845_ VGND VPWR VGND VPWR _07968_ keymem.key_mem\[9\]\[68\] _08377_ _08379_ _08380_
+ _07896_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_185_201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_154_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18352_ VPWR VGND VGND VPWR _04248_ _04249_ _04190_ sky130_fd_sc_hd__nor2_2
X_15564_ VGND VPWR _11023_ keymem.prev_key0_reg\[45\] keymem.prev_key0_reg\[77\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
X_12776_ VGND VPWR VGND VPWR _07547_ keymem.key_mem\[2\]\[61\] _08315_ _08317_ _08318_
+ _07662_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_201_588 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_115_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17303_ VPWR VGND VGND VPWR _11456_ _03399_ key[216] sky130_fd_sc_hd__nor2_2
X_14515_ VGND VPWR VGND VPWR _09982_ keymem.round_ctr_reg\[0\] _09984_ _09983_ sky130_fd_sc_hd__a21oi_2
X_11727_ VGND VPWR result[30] _07427_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15495_ VGND VPWR VPWR VGND _10955_ _10440_ _10953_ _10547_ _10954_ sky130_fd_sc_hd__o31a_2
X_18283_ VPWR VGND VGND VPWR _04185_ _04186_ _04077_ sky130_fd_sc_hd__nor2_2
XFILLER_0_126_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17234_ VPWR VGND VGND VPWR _03337_ key[209] _03077_ sky130_fd_sc_hd__nand2_2
X_14446_ VPWR VGND VGND VPWR _09329_ _09396_ _09915_ _09293_ _09623_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_83_298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11658_ VGND VPWR _00004_ _07392_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_9_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14377_ VPWR VGND VGND VPWR _09154_ _09847_ _09056_ sky130_fd_sc_hd__nor2_2
XFILLER_0_153_186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17165_ VGND VPWR VGND VPWR _03275_ _03274_ _10829_ _02708_ sky130_fd_sc_hd__o21a_2
XPHY_EDGE_ROW_167_2_Left_638 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_141_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_24_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16116_ VGND VPWR VGND VPWR _11569_ _11570_ _11464_ _11182_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_64_1537 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13328_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[116\] _07705_ keymem.key_mem\[4\]\[116\]
+ _07693_ _08815_ sky130_fd_sc_hd__a22o_2
XFILLER_0_12_538 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17096_ VPWR VGND VPWR VGND keymem.prev_key0_reg\[67\] _03213_ _09932_ _09985_ sky130_fd_sc_hd__or3b_2
XFILLER_0_126_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16047_ VGND VPWR VGND VPWR _11475_ _11501_ _11502_ _11300_ _11490_ sky130_fd_sc_hd__nor4_2
XFILLER_0_228_408 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13259_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[109\] _07724_ keymem.key_mem\[6\]\[109\]
+ _07565_ _08753_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_977 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_209_633 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_19_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19806_ VGND VPWR _00689_ _05312_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_97_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_986 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17998_ VPWR VGND VPWR VGND _03631_ _03930_ keymem.prev_key0_reg\[122\] _03788_ _00263_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_97_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19737_ VGND VPWR _00656_ _05276_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16949_ VGND VPWR VGND VPWR _02543_ _02542_ _02864_ _03080_ sky130_fd_sc_hd__a21o_2
XFILLER_0_205_850 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_206_Right_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_126_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19668_ VGND VPWR VPWR VGND _05091_ _05087_ keymem.key_mem\[12\]\[126\] _05238_ sky130_fd_sc_hd__mux2_2
XFILLER_0_232_680 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_133_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18619_ VPWR VGND _04488_ _04427_ enc_block.block_w0_reg\[3\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_137_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19599_ VPWR VGND keymem.key_mem\[12\]\[93\] _05202_ _05094_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_133_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21630_ VGND VPWR _01543_ _06282_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_176_267 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21561_ VGND VPWR VPWR VGND _06242_ _03592_ keymem.key_mem\[5\]\[116\] _06245_ sky130_fd_sc_hd__mux2_2
XFILLER_0_168_1318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_142_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_69_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_248_1320 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23300_ VGND VPWR _07182_ enc_block.round_key\[9\] _07181_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20512_ VGND VPWR _01020_ _05687_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_51_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24280_ VGND VPWR VPWR VGND clk _00773_ reset_n keymem.key_mem\[10\]\[17\] sky130_fd_sc_hd__dfrtp_2
X_21492_ VGND VPWR _01479_ _06208_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_69_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_490 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23231_ VPWR VGND _07119_ enc_block.block_w2_reg\[7\] enc_block.block_w2_reg\[2\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_215_Right_84 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20443_ VGND VPWR _00988_ _05650_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_31_814 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_259_500 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_144_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_696 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23162_ VGND VPWR VPWR VGND _07054_ _07065_ keymem.prev_key1_reg\[115\] _07066_ sky130_fd_sc_hd__mux2_2
XFILLER_0_67_1194 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20374_ VGND VPWR _05614_ _05533_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_109_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_144_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22113_ VGND VPWR VPWR VGND _06538_ _05069_ keymem.key_mem\[3\]\[117\] _06540_ sky130_fd_sc_hd__mux2_2
XFILLER_0_2_270 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_105_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23093_ VGND VPWR VGND VPWR _03413_ _03411_ _03416_ _07022_ sky130_fd_sc_hd__a21o_2
XFILLER_0_140_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22044_ VGND VPWR VPWR VGND _06494_ _05006_ keymem.key_mem\[3\]\[84\] _06504_ sky130_fd_sc_hd__mux2_2
XFILLER_0_105_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_485 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_76_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_224_Right_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25803_ keymem.prev_key1_reg\[119\] clk _02296_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_215_647 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_177_1171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23995_ VGND VPWR VPWR VGND clk _00488_ reset_n keymem.key_mem\[13\]\[116\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_216_1308 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25734_ keymem.prev_key1_reg\[50\] clk _02227_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22946_ VGND VPWR VGND VPWR _06935_ _02827_ _06891_ _02837_ _06892_ sky130_fd_sc_hd__a211o_2
XFILLER_0_253_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1010 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22877_ VGND VPWR _06892_ _06883_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25665_ VGND VPWR VPWR VGND clk _02158_ reset_n keymem.key_mem\[0\]\[122\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_167_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12630_ VGND VPWR VGND VPWR _07912_ keymem.key_mem\[11\]\[47\] _08183_ _08185_ _08186_
+ _08069_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_17_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24616_ VGND VPWR VPWR VGND clk _01109_ reset_n keymem.key_mem\[8\]\[97\] sky130_fd_sc_hd__dfrtp_2
X_21828_ VGND VPWR VPWR VGND _06377_ _03580_ keymem.key_mem\[4\]\[114\] _06386_ sky130_fd_sc_hd__mux2_2
XFILLER_0_39_947 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25596_ VGND VPWR VPWR VGND clk _02089_ reset_n keymem.key_mem\[0\]\[53\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_211_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_112_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1106 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_52_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24547_ VGND VPWR VPWR VGND clk _01040_ reset_n keymem.key_mem\[8\]\[28\] sky130_fd_sc_hd__dfrtp_2
X_12561_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[40\] _07536_ _08123_ _08119_ enc_block.round_key\[40\]
+ sky130_fd_sc_hd__o22a_2
X_21759_ VGND VPWR VPWR VGND _06344_ _03339_ keymem.key_mem\[4\]\[81\] _06350_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14300_ VGND VPWR VGND VPWR _09335_ _09343_ _09418_ _09495_ _09770_ sky130_fd_sc_hd__o22a_2
XFILLER_0_108_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15280_ VGND VPWR VGND VPWR _10740_ _10739_ _10743_ _10742_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_266_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24478_ VGND VPWR VPWR VGND clk _00971_ reset_n keymem.key_mem\[9\]\[87\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_237_Right_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12492_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[34\] _07924_ keymem.key_mem\[10\]\[34\]
+ _07562_ _08061_ sky130_fd_sc_hd__a22o_2
XFILLER_0_87_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14231_ VGND VPWR VGND VPWR _09702_ _09124_ _09646_ _09071_ _09040_ sky130_fd_sc_hd__a211o_2
X_23429_ VPWR VGND _07297_ _07167_ enc_block.block_w0_reg\[22\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_266_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14162_ VGND VPWR VGND VPWR _09631_ _09630_ _09632_ _09633_ sky130_fd_sc_hd__a21o_2
XFILLER_0_22_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13113_ VGND VPWR VGND VPWR _08622_ _08150_ keymem.key_mem\[3\]\[94\] _08619_ _08621_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_21_368 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14093_ VGND VPWR _09564_ _09563_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18970_ VPWR VGND VPWR VGND _04803_ block[54] _04744_ enc_block.block_w3_reg\[22\]
+ _04798_ _04804_ sky130_fd_sc_hd__a221o_2
XFILLER_0_81_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1036 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17921_ VGND VPWR _00238_ _03878_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13044_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[88\] _07652_ keymem.key_mem\[2\]\[88\]
+ _08116_ _08559_ sky130_fd_sc_hd__a22o_2
XFILLER_0_197_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17852_ VGND VPWR VGND VPWR _03289_ keymem.prev_key1_reg\[76\] _03831_ _03818_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_245_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_94_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16803_ VGND VPWR _02947_ _09517_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_227_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17783_ VGND VPWR VPWR VGND _03777_ _03783_ keymem.prev_key0_reg\[54\] _03784_ sky130_fd_sc_hd__mux2_2
X_14995_ VGND VPWR _10459_ _10458_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_238_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19522_ VGND VPWR VGND VPWR _05161_ keymem.key_mem_we _03109_ _05135_ _00556_ sky130_fd_sc_hd__a31o_2
XFILLER_0_221_606 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16734_ VGND VPWR VPWR VGND _02884_ keymem.key_mem\[14\]\[33\] _02883_ _02885_ sky130_fd_sc_hd__mux2_2
X_13946_ VGND VPWR _09418_ _09417_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_72_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_274 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_233_499 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_220_127 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_134_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19453_ VGND VPWR VGND VPWR _05124_ keymem.key_mem_we _02689_ _05121_ _00524_ sky130_fd_sc_hd__a31o_2
XFILLER_0_220_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_198_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16665_ VGND VPWR VGND VPWR _02586_ keymem.rcon_logic.tmp_rcon\[7\] _02819_ _02572_
+ sky130_fd_sc_hd__nand3_2
X_13877_ VGND VPWR _09349_ _09348_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18404_ VPWR VGND _04295_ _04127_ enc_block.block_w3_reg\[7\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15616_ VGND VPWR VGND VPWR _10481_ _10545_ _10504_ _10602_ _11074_ sky130_fd_sc_hd__o22a_2
XFILLER_0_57_722 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_134_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12828_ VPWR VGND VPWR VGND _08364_ keymem.key_mem\[9\]\[66\] _07919_ keymem.key_mem\[2\]\[66\]
+ _07647_ _08365_ sky130_fd_sc_hd__a221o_2
X_19384_ VGND VPWR VPWR VGND _05067_ _05083_ keymem.key_mem\[13\]\[124\] _05084_ sky130_fd_sc_hd__mux2_2
X_16596_ VGND VPWR _02753_ _02750_ _02752_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18335_ VPWR VGND VPWR VGND _04233_ _04189_ _04231_ enc_block.block_w0_reg\[23\]
+ _04097_ _00297_ sky130_fd_sc_hd__a221o_2
XFILLER_0_267_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15547_ VGND VPWR VGND VPWR _10480_ _10510_ _10563_ _10566_ _11006_ sky130_fd_sc_hd__o22a_2
XFILLER_0_210_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12759_ VPWR VGND VPWR VGND _08302_ keymem.key_mem\[5\]\[59\] _07683_ keymem.key_mem\[12\]\[59\]
+ _07621_ _08303_ sky130_fd_sc_hd__a221o_2
XFILLER_0_56_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18266_ VPWR VGND VPWR VGND _04170_ _04040_ _04168_ enc_block.block_w0_reg\[17\]
+ _04097_ _00291_ sky130_fd_sc_hd__a221o_2
X_15478_ VPWR VGND VPWR VGND _10938_ _10527_ _10618_ sky130_fd_sc_hd__or2_2
XFILLER_0_112_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_47_1009 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17217_ VGND VPWR _03322_ _03321_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14429_ VPWR VGND VPWR VGND _09472_ _09410_ _09478_ _09373_ _09898_ sky130_fd_sc_hd__or4_2
XFILLER_0_245_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18197_ VPWR VGND VGND VPWR _04107_ _04108_ _04041_ sky130_fd_sc_hd__nor2_2
XFILLER_0_126_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_181_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17148_ VGND VPWR VPWR VGND _03185_ keymem.key_mem\[14\]\[72\] _03259_ _03260_ sky130_fd_sc_hd__mux2_2
XFILLER_0_64_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17079_ VGND VPWR VGND VPWR _03197_ _03196_ _10386_ _03198_ sky130_fd_sc_hd__a21o_2
XFILLER_0_0_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20090_ VGND VPWR _00822_ _05463_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_224_411 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_174_1333 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22800_ VGND VPWR _06858_ _06779_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_27_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23780_ VPWR VGND VPWR VGND enc_block.ready reset_n _00273_ clk sky130_fd_sc_hd__dfstp_2
X_20992_ VGND VPWR _01244_ _05943_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_211_127 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22731_ VGND VPWR _02096_ _06830_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_211_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25450_ VGND VPWR VPWR VGND clk _01943_ reset_n keymem.key_mem\[1\]\[35\] sky130_fd_sc_hd__dfrtp_2
X_22662_ VGND VPWR _02055_ _06802_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_149_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1396 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_48_744 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24401_ VGND VPWR VPWR VGND clk _00894_ reset_n keymem.key_mem\[9\]\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_164_204 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21613_ VGND VPWR VGND VPWR _06259_ _10913_ _01535_ _06273_ sky130_fd_sc_hd__a21oi_2
X_25381_ VGND VPWR VPWR VGND clk _01874_ reset_n keymem.key_mem\[2\]\[94\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_34_1182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22593_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[105\] _06775_ _06774_ _05043_ _02013_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_1_1401 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_405 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_63_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24332_ VGND VPWR VPWR VGND clk _00825_ reset_n keymem.key_mem\[10\]\[69\] sky130_fd_sc_hd__dfrtp_2
X_21544_ VGND VPWR VPWR VGND _06231_ _03543_ keymem.key_mem\[5\]\[108\] _06236_ sky130_fd_sc_hd__mux2_2
XFILLER_0_7_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24263_ VGND VPWR VPWR VGND clk _00756_ reset_n keymem.key_mem\[10\]\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_105_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21475_ VPWR VGND VGND VPWR _06200_ keymem.key_mem\[5\]\[75\] _06114_ sky130_fd_sc_hd__nand2_2
XFILLER_0_16_674 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23214_ VPWR VGND VPWR VGND _07103_ block[1] _03958_ enc_block.block_w2_reg\[1\]
+ _03953_ _07104_ sky130_fd_sc_hd__a221o_2
X_20426_ VGND VPWR _00980_ _05641_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_244_1058 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24194_ VGND VPWR VPWR VGND clk _00687_ reset_n keymem.key_mem\[11\]\[59\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_30_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23145_ VGND VPWR VGND VPWR _07056_ _03540_ _06890_ _06924_ _03542_ sky130_fd_sc_hd__a211o_2
X_20357_ VGND VPWR _00947_ _05605_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_3_590 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_179_1211 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23076_ VGND VPWR VGND VPWR _03738_ key[210] _07013_ _03051_ sky130_fd_sc_hd__a21oi_2
X_20288_ VGND VPWR _05569_ _05534_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22027_ VGND VPWR VPWR VGND _06494_ _04992_ keymem.key_mem\[3\]\[76\] _06495_ sky130_fd_sc_hd__mux2_2
XFILLER_0_179_1255 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_255_1121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_76_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13800_ VPWR VGND VPWR VGND _09271_ _08985_ _09270_ _09269_ enc_block.block_w2_reg\[31\]
+ _09272_ sky130_fd_sc_hd__a221o_2
X_14780_ VGND VPWR VGND VPWR _09354_ _09474_ _09358_ _09443_ _10246_ sky130_fd_sc_hd__o22a_2
XFILLER_0_242_274 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11992_ VGND VPWR _07595_ _07594_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23978_ VGND VPWR VPWR VGND clk _00471_ reset_n keymem.key_mem\[13\]\[99\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_231_959 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_216_1149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_187_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13731_ VPWR VGND VPWR VGND _09031_ _09027_ _08971_ _08958_ _09203_ sky130_fd_sc_hd__or4_2
X_25717_ keymem.prev_key1_reg\[33\] clk _02210_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_97_143 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_192_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22929_ VGND VPWR VGND VPWR _02201_ _06923_ _06916_ keymem.prev_key1_reg\[24\] sky130_fd_sc_hd__o21a_2
XFILLER_0_196_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16450_ VPWR VGND VPWR VGND _02611_ _11570_ _11574_ sky130_fd_sc_hd__or2_2
XFILLER_0_42_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13662_ VGND VPWR _09134_ _09133_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25648_ VGND VPWR VPWR VGND clk _02141_ reset_n keymem.key_mem\[0\]\[105\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_116_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15401_ VGND VPWR VGND VPWR _10510_ _10411_ _10862_ _10459_ sky130_fd_sc_hd__a21oi_2
X_12613_ VPWR VGND VPWR VGND _08170_ keymem.key_mem\[5\]\[45\] _07597_ keymem.key_mem\[7\]\[45\]
+ _07610_ _08171_ sky130_fd_sc_hd__a221o_2
XFILLER_0_210_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13593_ VGND VPWR _09065_ _09064_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16381_ VPWR VGND VPWR VGND _02544_ keymem.prev_key0_reg\[21\] sky130_fd_sc_hd__inv_2
XFILLER_0_38_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25579_ VGND VPWR VPWR VGND clk _02072_ reset_n keymem.key_mem\[0\]\[36\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_155_248 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18120_ _04035_ _04037_ _04008_ _04036_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_15332_ VGND VPWR VGND VPWR _10441_ _10566_ _10521_ _10612_ _10794_ sky130_fd_sc_hd__o22a_2
XFILLER_0_26_427 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_87_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12544_ VPWR VGND VPWR VGND _08107_ keymem.key_mem\[3\]\[39\] _07844_ keymem.key_mem\[11\]\[39\]
+ _07781_ _08108_ sky130_fd_sc_hd__a221o_2
XFILLER_0_93_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18051_ VGND VPWR VGND VPWR _03972_ _09022_ _03973_ _03948_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_87_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15263_ VGND VPWR _10725_ _10628_ _10726_ _10490_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_48_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_268 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12475_ VGND VPWR enc_block.round_key\[32\] _08045_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_163_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_108_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17002_ VPWR VGND VPWR VGND _03128_ _10086_ _03125_ _03126_ _03127_ _10096_ sky130_fd_sc_hd__o311a_2
X_14214_ VGND VPWR VGND VPWR _09090_ _09684_ _09141_ _09127_ _09685_ sky130_fd_sc_hd__o22a_2
XFILLER_0_1_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15194_ VPWR VGND VPWR VGND _10658_ _10385_ sky130_fd_sc_hd__inv_2
XFILLER_0_227_1289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_806 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14145_ VGND VPWR VGND VPWR _09390_ _09340_ _09616_ _09378_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_240_1423 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_67_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18953_ VPWR VGND VGND VPWR _04778_ _04789_ _04201_ sky130_fd_sc_hd__nor2_2
X_14076_ VPWR VGND key[129] _09547_ _09511_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_226_709 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_24_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13027_ VGND VPWR VGND VPWR _07835_ keymem.key_mem\[13\]\[86\] _08541_ _08543_ _08544_
+ _08480_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_219_761 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17904_ VGND VPWR VGND VPWR _03792_ _02778_ _03727_ _03859_ _03867_ _03860_ sky130_fd_sc_hd__a2111o_2
X_18884_ VGND VPWR VGND VPWR _04725_ _03992_ _04726_ _00353_ sky130_fd_sc_hd__a21o_2
XFILLER_0_98_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17835_ VGND VPWR VPWR VGND _03814_ _03819_ keymem.prev_key0_reg\[70\] _03820_ sky130_fd_sc_hd__mux2_2
XFILLER_0_207_978 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_174_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_59_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_234_1205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_206_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17766_ VGND VPWR VPWR VGND _03763_ _03018_ keymem.prev_key0_reg\[47\] _03774_ sky130_fd_sc_hd__mux2_2
X_14978_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[12\] _08954_ _10442_ _08941_ _10417_
+ _10418_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_88_110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19505_ VGND VPWR _00548_ _05152_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16717_ VGND VPWR VPWR VGND _09523_ key[160] keymem.prev_key1_reg\[32\] _02869_ sky130_fd_sc_hd__mux2_2
X_13929_ VGND VPWR _09401_ _09400_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_57_1182 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17697_ VGND VPWR VPWR VGND _02947_ _03727_ _09534_ _03728_ sky130_fd_sc_hd__or3_2
XFILLER_0_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_88_176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19436_ VPWR VGND keymem.key_mem\[12\]\[17\] _05115_ _05102_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_9_605 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16648_ VGND VPWR VGND VPWR _02802_ _02801_ keymem.prev_key1_reg\[93\] _02803_ sky130_fd_sc_hd__a21o_2
XFILLER_0_57_541 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19367_ VGND VPWR _00490_ _05072_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_91_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16579_ VGND VPWR _02737_ keymem.prev_key1_reg\[26\] keymem.prev_key1_reg\[58\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_169_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18318_ _04216_ _04218_ _04215_ _04217_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_267_1058 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19298_ VGND VPWR VPWR VGND _05025_ _05024_ keymem.key_mem\[13\]\[96\] _05026_ sky130_fd_sc_hd__mux2_2
XFILLER_0_33_909 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_169_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_66_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18249_ VPWR VGND VPWR VGND _04155_ _04079_ _04153_ sky130_fd_sc_hd__or2_2
XFILLER_0_154_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_6_Right_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_199_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_199_79 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21260_ VGND VPWR _01370_ _06085_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_41_953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20211_ VGND VPWR _00880_ _05526_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_100_2_Left_571 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21191_ VGND VPWR _01337_ _06049_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_243_1091 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_106_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20142_ VGND VPWR _00847_ _05490_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_110_395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24950_ VGND VPWR VPWR VGND clk _01443_ reset_n keymem.key_mem\[5\]\[47\] sky130_fd_sc_hd__dfrtp_2
X_20073_ VGND VPWR _00814_ _05454_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_148_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23901_ VGND VPWR VPWR VGND clk _00394_ reset_n keymem.key_mem\[13\]\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_256_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24881_ VGND VPWR VPWR VGND clk _01374_ reset_n keymem.key_mem\[6\]\[106\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_1_Left_418 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23832_ VGND VPWR VPWR VGND clk _00325_ reset_n enc_block.block_w1_reg\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_256_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1174 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_217_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23763_ keymem.prev_key0_reg\[119\] clk _00260_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20975_ VGND VPWR VPWR VGND _05934_ _05024_ keymem.key_mem\[7\]\[96\] _05935_ sky130_fd_sc_hd__mux2_2
XFILLER_0_67_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_778 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25502_ VGND VPWR VPWR VGND clk _01995_ reset_n keymem.key_mem\[1\]\[87\] sky130_fd_sc_hd__dfrtp_2
X_22714_ VGND VPWR VPWR VGND _06822_ keymem.key_mem\[0\]\[51\] _03068_ _06823_ sky130_fd_sc_hd__mux2_2
XFILLER_0_113_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23694_ keymem.prev_key0_reg\[50\] clk _00191_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_67_349 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_250_1084 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22645_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[11\] _06790_ _06789_ _04894_ _02047_
+ sky130_fd_sc_hd__a22o_2
X_25433_ VGND VPWR VPWR VGND clk _01926_ reset_n keymem.key_mem\[1\]\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_187_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25364_ VGND VPWR VPWR VGND clk _01857_ reset_n keymem.key_mem\[2\]\[77\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_192_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_75_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22576_ VGND VPWR _02000_ _06771_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_148_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_84_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24315_ VGND VPWR VPWR VGND clk _00808_ reset_n keymem.key_mem\[10\]\[52\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_267_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21527_ VGND VPWR VPWR VGND _06220_ _03492_ keymem.key_mem\[5\]\[100\] _06227_ sky130_fd_sc_hd__mux2_2
X_25295_ VGND VPWR VPWR VGND clk _01788_ reset_n keymem.key_mem\[2\]\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_228_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24246_ VGND VPWR VPWR VGND clk _00739_ reset_n keymem.key_mem\[11\]\[111\] sky130_fd_sc_hd__dfrtp_2
X_12260_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[14\] _07536_ _07848_ _07837_ enc_block.round_key\[14\]
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_259_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21458_ VGND VPWR VPWR VGND _06184_ _03216_ keymem.key_mem\[5\]\[67\] _06191_ sky130_fd_sc_hd__mux2_2
XFILLER_0_224_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20409_ VGND VPWR _00972_ _05632_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24177_ VGND VPWR VPWR VGND clk _00670_ reset_n keymem.key_mem\[11\]\[42\] sky130_fd_sc_hd__dfrtp_2
X_12191_ VPWR VGND VPWR VGND _07783_ keymem.key_mem\[5\]\[10\] _07780_ keymem.key_mem\[3\]\[10\]
+ _07778_ _07784_ sky130_fd_sc_hd__a221o_2
XFILLER_0_160_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21389_ VGND VPWR VPWR VGND _06151_ _02893_ keymem.key_mem\[5\]\[34\] _06155_ sky130_fd_sc_hd__mux2_2
XFILLER_0_43_1226 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23128_ VGND VPWR _02279_ _07044_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_124_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15950_ VPWR VGND VPWR VGND _11394_ _11405_ _11401_ _11388_ _11406_ sky130_fd_sc_hd__or4_2
X_23059_ VGND VPWR VPWR VGND _06992_ _07002_ keymem.prev_key1_reg\[75\] _07003_ sky130_fd_sc_hd__mux2_2
X_14901_ VGND VPWR _10366_ _09987_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15881_ VGND VPWR VGND VPWR _11336_ _11205_ _11337_ _11314_ sky130_fd_sc_hd__a21oi_2
X_17620_ VGND VPWR _03675_ _03674_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14832_ VPWR VGND VPWR VGND _09328_ _09476_ _09339_ _09338_ _10297_ sky130_fd_sc_hd__or4_2
XFILLER_0_235_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_403 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_192_1263 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_235_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17551_ VPWR VGND VGND VPWR _03615_ _03240_ _02672_ sky130_fd_sc_hd__nand2_2
XFILLER_0_8_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14763_ VPWR VGND VGND VPWR _09075_ _10222_ _10228_ _10229_ sky130_fd_sc_hd__nor3_2
XPHY_EDGE_ROW_176_2_Left_647 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_153_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11975_ VGND VPWR _07578_ _07577_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16502_ VGND VPWR VPWR VGND _02662_ keymem.key_mem\[14\]\[23\] _02661_ _02663_ sky130_fd_sc_hd__mux2_2
X_13714_ VPWR VGND VGND VPWR _09186_ _09184_ _09185_ sky130_fd_sc_hd__nand2_2
X_17482_ VGND VPWR VPWR VGND _03534_ keymem.key_mem\[14\]\[110\] _03555_ _03556_ sky130_fd_sc_hd__mux2_2
XFILLER_0_39_530 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14694_ VGND VPWR VGND VPWR _09221_ _09110_ _09149_ _09160_ _10161_ sky130_fd_sc_hd__o22a_2
XFILLER_0_170_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19221_ VGND VPWR _00438_ _04978_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_224_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16433_ VGND VPWR VGND VPWR _09517_ _02593_ _02591_ _02592_ _02595_ sky130_fd_sc_hd__a31o_2
XFILLER_0_27_703 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13645_ VGND VPWR VGND VPWR _09107_ _09113_ _09116_ _09114_ _09117_ sky130_fd_sc_hd__o22a_2
XFILLER_0_195_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_736 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19152_ VGND VPWR VPWR VGND _04928_ _04935_ keymem.key_mem\[13\]\[40\] _04936_ sky130_fd_sc_hd__mux2_2
XFILLER_0_27_747 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16364_ _11409_ _02527_ _11258_ _11417_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_54_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13576_ VGND VPWR VPWR VGND _09042_ _09040_ _09048_ _09047_ _09046_ sky130_fd_sc_hd__o211a_2
XFILLER_0_183_387 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18103_ VPWR VGND _04021_ enc_block.block_w0_reg\[31\] enc_block.block_w0_reg\[27\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_59_Right_59 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15315_ _10487_ _10777_ _10764_ _10765_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_12527_ VPWR VGND VPWR VGND _08092_ keymem.key_mem\[9\]\[37\] _07672_ keymem.key_mem\[8\]\[37\]
+ _07541_ _08093_ sky130_fd_sc_hd__a221o_2
X_19083_ VGND VPWR _00383_ _04895_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_41_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16295_ VGND VPWR VGND VPWR _02458_ _02430_ _07386_ _02459_ sky130_fd_sc_hd__a21o_2
X_18034_ VPWR VGND VGND VPWR _03955_ _03956_ _03947_ sky130_fd_sc_hd__nor2_2
X_15246_ VPWR VGND VGND VPWR _10476_ _10709_ _10608_ sky130_fd_sc_hd__nor2_2
XFILLER_0_23_942 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_23_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12458_ VPWR VGND VPWR VGND _08029_ keymem.key_mem\[10\]\[31\] _07561_ keymem.key_mem\[12\]\[31\]
+ _07578_ _08030_ sky130_fd_sc_hd__a221o_2
XFILLER_0_169_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15177_ VPWR VGND VGND VPWR _10511_ _10639_ _10641_ _10547_ _10635_ sky130_fd_sc_hd__o22ai_2
X_12389_ VGND VPWR VGND VPWR _07542_ keymem.key_mem\[8\]\[25\] _07964_ _07966_ _07967_
+ _07663_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_61_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14128_ VPWR VGND VGND VPWR _09410_ _09599_ _09268_ sky130_fd_sc_hd__nor2_2
XFILLER_0_240_1253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19985_ VGND VPWR _00772_ _05408_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_185_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_377 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18936_ VGND VPWR _04773_ _04711_ _04772_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_14059_ VPWR VGND VGND VPWR _09531_ _09529_ _09530_ sky130_fd_sc_hd__nand2_2
XFILLER_0_94_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18867_ VPWR VGND _04711_ enc_block.block_w0_reg\[15\] enc_block.block_w0_reg\[11\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_59_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_222_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17818_ VGND VPWR _00206_ _03807_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_265_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18798_ VPWR VGND VPWR VGND _04649_ _04646_ _04648_ sky130_fd_sc_hd__or2_2
XFILLER_0_94_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17749_ VGND VPWR VPWR VGND _03763_ _02951_ keymem.prev_key0_reg\[40\] _03764_ sky130_fd_sc_hd__mux2_2
XFILLER_0_171_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20760_ VGND VPWR VPWR VGND _05679_ _03668_ keymem.key_mem\[8\]\[127\] _05817_ sky130_fd_sc_hd__mux2_2
XFILLER_0_58_850 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_72_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_134_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19419_ VPWR VGND keymem.key_mem\[12\]\[9\] _05106_ _05102_ VPWR VGND sky130_fd_sc_hd__and2_2
X_20691_ VGND VPWR VPWR VGND _05772_ _03452_ keymem.key_mem\[8\]\[94\] _05781_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_1141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22430_ VGND VPWR VPWR VGND _06702_ keymem.key_mem\[1\]\[9\] _10747_ _06709_ sky130_fd_sc_hd__mux2_2
XFILLER_0_174_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_18_769 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_94_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22361_ VGND VPWR _01885_ _06671_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24100_ VGND VPWR VPWR VGND clk _00593_ reset_n keymem.key_mem\[12\]\[93\] sky130_fd_sc_hd__dfrtp_2
X_21312_ VGND VPWR _01395_ _06112_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25080_ VGND VPWR VPWR VGND clk _01573_ reset_n keymem.key_mem\[4\]\[49\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_182_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22292_ VGND VPWR _01852_ _06635_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_5_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_206_1126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24031_ VGND VPWR VPWR VGND clk _00524_ reset_n keymem.key_mem\[12\]\[24\] sky130_fd_sc_hd__dfrtp_2
X_21243_ VGND VPWR VPWR VGND _06076_ _03452_ keymem.key_mem\[6\]\[94\] _06077_ sky130_fd_sc_hd__mux2_2
XFILLER_0_182_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21174_ VGND VPWR VPWR VGND _06040_ _03161_ keymem.key_mem\[6\]\[61\] _06041_ sky130_fd_sc_hd__mux2_2
XFILLER_0_256_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_141_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20125_ VGND VPWR _00839_ _05481_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_217_517 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_102_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_77_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20056_ VGND VPWR _00806_ _05445_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24933_ VGND VPWR VPWR VGND clk _01426_ reset_n keymem.key_mem\[5\]\[30\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24864_ VGND VPWR VPWR VGND clk _01357_ reset_n keymem.key_mem\[6\]\[89\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_225_583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_252_1124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_193_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23815_ VGND VPWR VPWR VGND clk _00308_ reset_n enc_block.block_w1_reg\[0\] sky130_fd_sc_hd__dfrtp_2
X_24795_ VGND VPWR VPWR VGND clk _01288_ reset_n keymem.key_mem\[6\]\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11760_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[15\] dec_new_block\[47\]
+ _07444_ sky130_fd_sc_hd__mux2_2
XFILLER_0_90_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23746_ keymem.prev_key0_reg\[102\] clk _00243_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20958_ VGND VPWR VPWR VGND _05912_ _05013_ keymem.key_mem\[7\]\[88\] _05926_ sky130_fd_sc_hd__mux2_2
XFILLER_0_261_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11691_ VGND VPWR result[12] _07409_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_49_872 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23677_ keymem.prev_key0_reg\[33\] clk _00174_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20889_ VGND VPWR _01195_ _05889_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_230_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_187_1332 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13430_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[126\] _07924_ keymem.key_mem\[11\]\[126\]
+ _08090_ _08907_ sky130_fd_sc_hd__a22o_2
X_25416_ VGND VPWR VPWR VGND clk _01909_ reset_n keymem.key_mem\[1\]\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_36_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_125_207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22628_ VGND VPWR _06784_ _06778_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_64_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1376 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_49_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13361_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[119\] _07651_ keymem.key_mem\[6\]\[119\]
+ _07656_ _08845_ sky130_fd_sc_hd__a22o_2
XFILLER_0_63_363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25347_ VGND VPWR VPWR VGND clk _01840_ reset_n keymem.key_mem\[2\]\[60\] sky130_fd_sc_hd__dfrtp_2
X_22559_ VGND VPWR _01990_ _06764_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_64_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15100_ VPWR VGND VGND VPWR _10520_ _10564_ _10563_ sky130_fd_sc_hd__nor2_2
XFILLER_0_49_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12312_ VGND VPWR _07896_ _07662_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16080_ VGND VPWR _11534_ _11458_ _11535_ _11533_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_13292_ VPWR VGND VPWR VGND _08782_ keymem.key_mem\[13\]\[112\] _08125_ keymem.key_mem\[2\]\[112\]
+ _07647_ _08783_ sky130_fd_sc_hd__a221o_2
X_25278_ VGND VPWR VPWR VGND clk _01771_ reset_n keymem.key_mem\[3\]\[119\] sky130_fd_sc_hd__dfrtp_2
X_15031_ VGND VPWR _10495_ _10494_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12243_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[14\] _07609_ keymem.key_mem\[2\]\[14\]
+ _07546_ _07832_ sky130_fd_sc_hd__a22o_2
XFILLER_0_161_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24229_ VGND VPWR VPWR VGND clk _00722_ reset_n keymem.key_mem\[11\]\[94\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_934 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12174_ VPWR VGND VPWR VGND _07767_ keymem.key_mem\[14\]\[9\] _07632_ keymem.key_mem\[11\]\[9\]
+ _07631_ _07768_ sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_170_2_Right_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19770_ VGND VPWR VPWR VGND _05292_ keymem.key_mem\[11\]\[44\] _02998_ _05294_ sky130_fd_sc_hd__mux2_2
X_16982_ VGND VPWR VPWR VGND _03084_ keymem.key_mem\[14\]\[56\] _03109_ _03110_ sky130_fd_sc_hd__mux2_2
XFILLER_0_159_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18721_ VPWR VGND VPWR VGND _04579_ _04434_ _04577_ sky130_fd_sc_hd__or2_2
X_15933_ VPWR VGND VGND VPWR _11286_ _11389_ _11376_ sky130_fd_sc_hd__nor2_2
XFILLER_0_218_1008 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18652_ VPWR VGND VGND VPWR _04517_ _04518_ _04478_ sky130_fd_sc_hd__nor2_2
X_15864_ VGND VPWR _11320_ _11319_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17603_ VPWR VGND VPWR VGND _03660_ _03657_ _03656_ key[254] _08929_ _03661_ sky130_fd_sc_hd__a221o_2
XFILLER_0_235_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14815_ VGND VPWR _10281_ _07378_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18583_ _04454_ _04456_ _04294_ _04455_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_15795_ VPWR VGND VPWR VGND _11206_ _11202_ _11197_ _11187_ _11251_ sky130_fd_sc_hd__or4_2
XFILLER_0_231_1219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17534_ VGND VPWR VPWR VGND _03593_ keymem.key_mem\[14\]\[117\] _03600_ _03601_ sky130_fd_sc_hd__mux2_2
X_14746_ VGND VPWR VPWR VGND _09108_ _09157_ _09228_ _10212_ sky130_fd_sc_hd__or3_2
XFILLER_0_59_647 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11958_ VGND VPWR _07561_ _07560_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_54_1174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17465_ VPWR VGND VGND VPWR _03541_ key[236] _10967_ sky130_fd_sc_hd__nand2_2
X_14677_ VPWR VGND VGND VPWR _10144_ _09732_ _10143_ sky130_fd_sc_hd__nand2_2
X_11889_ VGND VPWR result[111] _07508_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_15_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19204_ VPWR VGND keymem.key_mem\[13\]\[59\] _04969_ _04961_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16416_ VPWR VGND VPWR VGND _02451_ _02577_ _02576_ _02450_ _02578_ sky130_fd_sc_hd__or4_2
X_13628_ VGND VPWR _09100_ _09099_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_156_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17396_ VGND VPWR _00110_ _03481_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19135_ VPWR VGND keymem.key_mem\[13\]\[34\] _04925_ _04915_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_264_1017 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16347_ VGND VPWR VGND VPWR _11352_ _11305_ _11238_ _11361_ _02510_ sky130_fd_sc_hd__o22a_2
XFILLER_0_55_886 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_109_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13559_ VGND VPWR _09031_ _09030_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_55_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_67_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19066_ VGND VPWR VGND VPWR _04885_ keymem.key_mem_we _10099_ _04878_ _00376_ sky130_fd_sc_hd__a31o_2
XFILLER_0_14_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16278_ VGND VPWR VGND VPWR _02441_ _11323_ _11230_ _11291_ _02442_ sky130_fd_sc_hd__a31o_2
XFILLER_0_42_569 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_207_1446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_2_633 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18017_ VGND VPWR VGND VPWR _03941_ enc_block.round\[1\] _03943_ _00000_ sky130_fd_sc_hd__a21oi_2
X_15229_ VPWR VGND VPWR VGND _10689_ _10691_ _10690_ _10688_ _10692_ sky130_fd_sc_hd__or4_2
XFILLER_0_207_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_433 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_201_1001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_239_664 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_11_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19968_ VGND VPWR VPWR VGND _05389_ _10747_ keymem.key_mem\[10\]\[9\] _05399_ sky130_fd_sc_hd__mux2_2
XFILLER_0_96_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18919_ VPWR VGND VGND VPWR _04757_ _04758_ _04478_ sky130_fd_sc_hd__nor2_2
XFILLER_0_138_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19899_ VGND VPWR _05361_ _05242_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_59_1030 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_207_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21930_ VPWR VGND keymem.key_mem\[3\]\[31\] _06443_ _06439_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_218_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21861_ VPWR VGND VGND VPWR _06405_ _08933_ _05241_ sky130_fd_sc_hd__nand2_2
X_23600_ VGND VPWR VPWR VGND clk _00101_ reset_n keymem.key_mem\[14\]\[89\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_239_Left_506 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20812_ VPWR VGND keymem.key_mem\[7\]\[20\] _05848_ _05844_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_136_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21792_ VGND VPWR _01620_ _06367_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24580_ VGND VPWR VPWR VGND clk _01073_ reset_n keymem.key_mem\[8\]\[61\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_72_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20743_ VGND VPWR _01130_ _05808_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23531_ VGND VPWR VPWR VGND clk _00032_ reset_n keymem.key_mem\[14\]\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_522 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23462_ VGND VPWR _07326_ _04256_ _02331_ _07096_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_20674_ VGND VPWR _05772_ _05675_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_107_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25201_ VGND VPWR VPWR VGND clk _01694_ reset_n keymem.key_mem\[3\]\[42\] sky130_fd_sc_hd__dfrtp_2
X_22413_ VGND VPWR VPWR VGND _06696_ keymem.key_mem\[1\]\[2\] _09862_ _06699_ sky130_fd_sc_hd__mux2_2
X_23393_ VGND VPWR _07265_ _07204_ _07264_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22344_ VGND VPWR _01877_ _06662_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25132_ VGND VPWR VPWR VGND clk _01625_ reset_n keymem.key_mem\[4\]\[101\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_225_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_248_Left_515 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25063_ VGND VPWR VPWR VGND clk _01556_ reset_n keymem.key_mem\[4\]\[32\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22275_ VGND VPWR _01844_ _06626_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_143_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24014_ VGND VPWR VPWR VGND clk _00507_ reset_n keymem.key_mem\[12\]\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_104_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21226_ VGND VPWR VPWR VGND _06065_ _03383_ keymem.key_mem\[6\]\[86\] _06068_ sky130_fd_sc_hd__mux2_2
XFILLER_0_130_276 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_143_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21157_ VGND VPWR VPWR VGND _06029_ _03082_ keymem.key_mem\[6\]\[53\] _06032_ sky130_fd_sc_hd__mux2_2
XFILLER_0_244_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20108_ VPWR VGND VGND VPWR _05473_ keymem.key_mem\[10\]\[75\] _05402_ sky130_fd_sc_hd__nand2_2
X_21088_ VGND VPWR _01288_ _05995_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12930_ VGND VPWR VGND VPWR _08457_ _08050_ keymem.key_mem\[7\]\[76\] _08454_ _08456_
+ sky130_fd_sc_hd__a211o_2
X_20039_ VGND VPWR VPWR VGND _05435_ _02972_ keymem.key_mem\[10\]\[42\] _05437_ sky130_fd_sc_hd__mux2_2
X_24916_ VGND VPWR VPWR VGND clk _01409_ reset_n keymem.key_mem\[5\]\[13\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_257_Left_524 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_87_219 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12861_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[69\] _08259_ _08394_ _08389_ _08395_
+ sky130_fd_sc_hd__o22a_2
X_24847_ VGND VPWR VPWR VGND clk _01340_ reset_n keymem.key_mem\[6\]\[72\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14600_ VPWR VGND VGND VPWR _09386_ _10068_ _09312_ sky130_fd_sc_hd__nor2_2
XFILLER_0_154_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11812_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[9\] dec_new_block\[73\]
+ _07470_ sky130_fd_sc_hd__mux2_2
X_15580_ VPWR VGND VPWR VGND _11038_ _10085_ _11029_ key[141] _09544_ _11039_ sky130_fd_sc_hd__a221o_2
X_12792_ VGND VPWR enc_block.round_key\[62\] _08332_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24778_ VGND VPWR VPWR VGND clk _01271_ reset_n keymem.key_mem\[6\]\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_90_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_189_1405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14531_ VGND VPWR VGND VPWR _09145_ _09684_ _09999_ _09132_ sky130_fd_sc_hd__a21oi_2
X_11743_ VGND VPWR result[38] _07435_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23729_ keymem.prev_key0_reg\[85\] clk _00226_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_3_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17250_ VGND VPWR VGND VPWR _03351_ _09513_ _10732_ key[83] sky130_fd_sc_hd__o21a_2
XFILLER_0_138_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14462_ VGND VPWR _09931_ _09512_ VPWR VGND sky130_fd_sc_hd__buf_1
X_11674_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[4\] dec_new_block\[4\]
+ _07401_ sky130_fd_sc_hd__mux2_2
X_16201_ VGND VPWR VGND VPWR _11218_ _11250_ _02366_ _11404_ sky130_fd_sc_hd__a21oi_2
X_13413_ VGND VPWR VGND VPWR _07842_ keymem.key_mem\[9\]\[124\] _08887_ _08889_ _08892_
+ _08891_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_3_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17181_ VPWR VGND VGND VPWR _03289_ key[204] _10967_ sky130_fd_sc_hd__nand2_2
XFILLER_0_37_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14393_ VGND VPWR _09863_ _09540_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16132_ VGND VPWR VGND VPWR _11400_ _11367_ _11239_ _11386_ _11586_ sky130_fd_sc_hd__o22a_2
XPHY_EDGE_ROW_266_Left_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13344_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[117\] _08714_ _08829_ _08825_ _08830_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_84_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16063_ VGND VPWR VGND VPWR _11204_ _11295_ _11250_ _11464_ _11518_ sky130_fd_sc_hd__o22a_2
XFILLER_0_11_219 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13275_ VGND VPWR VGND VPWR _08768_ _07580_ keymem.key_mem\[12\]\[110\] _08765_ _08767_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_62_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_161_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15014_ VPWR VGND VGND VPWR _10478_ _10463_ _10477_ sky130_fd_sc_hd__nand2_2
XFILLER_0_122_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12226_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[12\] _07629_ keymem.key_mem\[2\]\[12\]
+ _07816_ _07817_ sky130_fd_sc_hd__a22o_2
XFILLER_0_20_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_255_409 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_161_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19822_ VGND VPWR VPWR VGND _05314_ keymem.key_mem\[11\]\[69\] _03235_ _05321_ sky130_fd_sc_hd__mux2_2
X_12157_ VGND VPWR _07752_ _07539_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_23_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_75_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_171_2_Right_243 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16965_ VGND VPWR VGND VPWR _03094_ _10328_ _02877_ key[55] sky130_fd_sc_hd__o21a_2
X_19753_ VGND VPWR VPWR VGND _05281_ keymem.key_mem\[11\]\[36\] _02913_ _05285_ sky130_fd_sc_hd__mux2_2
X_12088_ VPWR VGND VPWR VGND _07686_ keymem.key_mem\[14\]\[4\] _07685_ keymem.key_mem\[6\]\[4\]
+ _07639_ _07687_ sky130_fd_sc_hd__a221o_2
XFILLER_0_251_626 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15916_ VGND VPWR _11372_ _11334_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18704_ VPWR VGND VPWR VGND _04564_ _04353_ _04562_ sky130_fd_sc_hd__or2_2
X_19684_ VGND VPWR VPWR VGND _05247_ keymem.key_mem\[11\]\[3\] _09992_ _05249_ sky130_fd_sc_hd__mux2_2
X_16896_ VGND VPWR VPWR VGND _09523_ key[176] keymem.prev_key1_reg\[48\] _03032_ sky130_fd_sc_hd__mux2_2
XFILLER_0_216_380 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18635_ VPWR VGND VGND VPWR _04380_ _04503_ _04201_ sky130_fd_sc_hd__nor2_2
XFILLER_0_78_208 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_188_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15847_ VGND VPWR _11303_ _11302_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_95_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_172_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_133_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_152_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18566_ VPWR VGND _04441_ _04440_ enc_block.round_key\[77\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_115_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15778_ VGND VPWR VPWR VGND _11173_ _11180_ _11233_ _11234_ sky130_fd_sc_hd__or3_2
XFILLER_0_24_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_133_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17517_ VGND VPWR VPWR VGND _03534_ keymem.key_mem\[14\]\[115\] _03585_ _03586_ sky130_fd_sc_hd__mux2_2
X_14729_ VGND VPWR _00017_ _10195_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18497_ VPWR VGND _04379_ _04378_ enc_block.round_key\[70\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_24_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17448_ VGND VPWR _00117_ _03526_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_131_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17379_ VGND VPWR _03467_ _09540_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_15_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_27_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19118_ VGND VPWR VGND VPWR _04914_ keymem.key_mem_we _02765_ _04908_ _00399_ sky130_fd_sc_hd__a31o_2
XFILLER_0_171_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_867 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20390_ VGND VPWR _00963_ _05622_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_160_1_Left_427 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_183_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19049_ VGND VPWR _04874_ _03949_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_242_1123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_144_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22060_ VPWR VGND keymem.key_mem\[3\]\[92\] _06512_ _06405_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_80_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_220_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21011_ VGND VPWR _01253_ _05953_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_57_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25750_ keymem.prev_key1_reg\[66\] clk _02243_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22962_ VPWR VGND VGND VPWR _06881_ _06945_ keymem.prev_key1_reg\[36\] sky130_fd_sc_hd__nor2_2
XFILLER_0_65_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24701_ VGND VPWR VPWR VGND clk _01194_ reset_n keymem.key_mem\[7\]\[54\] sky130_fd_sc_hd__dfrtp_2
X_21913_ VPWR VGND keymem.key_mem\[3\]\[23\] _06434_ _06427_ VPWR VGND sky130_fd_sc_hd__and2_2
X_25681_ VGND VPWR VPWR VGND clk _02174_ reset_n keymem.round_ctr_reg\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_190_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22893_ VGND VPWR VPWR VGND _06878_ _06901_ keymem.prev_key1_reg\[10\] _06902_ sky130_fd_sc_hd__mux2_2
XFILLER_0_151_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24632_ VGND VPWR VPWR VGND clk _01125_ reset_n keymem.key_mem\[8\]\[113\] sky130_fd_sc_hd__dfrtp_2
X_21844_ VGND VPWR _01645_ _06394_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_190_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_151_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24563_ VGND VPWR VPWR VGND clk _01056_ reset_n keymem.key_mem\[8\]\[44\] sky130_fd_sc_hd__dfrtp_2
X_21775_ VGND VPWR _01612_ _06358_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_231_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_194_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_80 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23514_ VGND VPWR VPWR VGND clk _00015_ reset_n keymem.key_mem\[14\]\[3\] sky130_fd_sc_hd__dfrtp_2
X_20726_ VGND VPWR _01122_ _05799_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_4_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24494_ VGND VPWR VPWR VGND clk _00987_ reset_n keymem.key_mem\[9\]\[103\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_875 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_247_1012 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23445_ VPWR VGND VPWR VGND _07311_ _03950_ _07310_ enc_block.block_w3_reg\[24\]
+ _07126_ _02329_ sky130_fd_sc_hd__a221o_2
X_20657_ VGND VPWR _01089_ _05763_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_18_385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_92_1_Left_359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23376_ VPWR VGND VGND VPWR _07250_ _07247_ _07249_ sky130_fd_sc_hd__nand2_2
X_20588_ VGND VPWR _01056_ _05727_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25115_ VGND VPWR VPWR VGND clk _01608_ reset_n keymem.key_mem\[4\]\[84\] sky130_fd_sc_hd__dfrtp_2
X_22327_ VGND VPWR _01869_ _06653_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_249_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13060_ VPWR VGND VPWR VGND _08573_ keymem.key_mem\[14\]\[89\] _07706_ keymem.key_mem\[9\]\[89\]
+ _07919_ _08574_ sky130_fd_sc_hd__a221o_2
X_22258_ VGND VPWR _01836_ _06617_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25046_ VGND VPWR VPWR VGND clk _01539_ reset_n keymem.key_mem\[4\]\[15\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_185_2_Left_656 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12011_ VGND VPWR _07613_ _07595_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21209_ VGND VPWR VPWR VGND _06052_ _03314_ keymem.key_mem\[6\]\[78\] _06059_ sky130_fd_sc_hd__mux2_2
X_22189_ VGND VPWR _01803_ _06581_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_44_1195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_217_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_79_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16750_ VPWR VGND _10366_ _02899_ _09985_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_245_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_233_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13962_ VGND VPWR _09434_ _09433_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_96_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_254_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_147 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15701_ VGND VPWR VPWR VGND _08927_ _11156_ key[144] _11157_ sky130_fd_sc_hd__mux2_2
X_12913_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[75\] _07843_ keymem.key_mem\[10\]\[75\]
+ _08193_ _08441_ sky130_fd_sc_hd__a22o_2
X_16681_ VGND VPWR VGND VPWR _02832_ _02831_ _02835_ _02833_ sky130_fd_sc_hd__a21oi_2
X_13893_ VPWR VGND VPWR VGND _09307_ _09308_ _09285_ _09338_ _09365_ sky130_fd_sc_hd__or4_2
X_18420_ VGND VPWR _04308_ enc_block.block_w1_reg\[24\] _04307_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15632_ VGND VPWR VPWR VGND _11072_ _11089_ _09240_ _11090_ sky130_fd_sc_hd__or3_2
X_12844_ VPWR VGND VPWR VGND _08378_ keymem.key_mem\[3\]\[68\] _08216_ keymem.key_mem\[8\]\[68\]
+ _07541_ _08379_ sky130_fd_sc_hd__a221o_2
XFILLER_0_154_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18351_ VGND VPWR VGND VPWR _09629_ _09589_ _04073_ _04248_ sky130_fd_sc_hd__a21o_2
XFILLER_0_61_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15563_ VGND VPWR VGND VPWR _11020_ _11019_ _10979_ _11022_ sky130_fd_sc_hd__a21o_2
XFILLER_0_90_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12775_ VPWR VGND VPWR VGND _08316_ keymem.key_mem\[14\]\[61\] _07632_ keymem.key_mem\[4\]\[61\]
+ _07692_ _08317_ sky130_fd_sc_hd__a221o_2
X_17302_ VGND VPWR VGND VPWR key[88] _08937_ _03397_ _03396_ _03398_ sky130_fd_sc_hd__o22a_2
X_14514_ _09883_ _09983_ _07386_ _09923_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_232_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18282_ VGND VPWR _04185_ _04182_ _04184_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_11726_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[30\] dec_new_block\[30\]
+ _07427_ sky130_fd_sc_hd__mux2_2
X_15494_ VGND VPWR VGND VPWR _10609_ _10583_ _10501_ _10867_ _10954_ sky130_fd_sc_hd__o22a_2
XFILLER_0_16_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_458 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_126_324 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17233_ VGND VPWR VGND VPWR _03336_ _03302_ _02927_ key[81] sky130_fd_sc_hd__o21a_2
XFILLER_0_86_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_335 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_232_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14445_ VGND VPWR VGND VPWR _09623_ _09486_ _09914_ _09311_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_193_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11657_ VGND VPWR VPWR VGND _07371_ aes_core_ctrl_reg\[0\] _07391_ _07392_ sky130_fd_sc_hd__mux2_2
X_17164_ VPWR VGND VGND VPWR _03274_ key[202] _10092_ sky130_fd_sc_hd__nand2_2
X_14376_ VPWR VGND VGND VPWR _09216_ _09174_ _09846_ _09100_ _09156_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_208_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16115_ _11291_ _11569_ _11395_ _11408_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_141_349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13327_ VGND VPWR VGND VPWR _08814_ _07877_ keymem.key_mem\[10\]\[116\] _08813_ _08020_
+ sky130_fd_sc_hd__a211o_2
X_17095_ VPWR VGND VGND VPWR _03212_ _10189_ _09985_ sky130_fd_sc_hd__nand2_2
XFILLER_0_10_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_78 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16046_ VGND VPWR VPWR VGND _11496_ _11500_ _11492_ _11501_ sky130_fd_sc_hd__or3_2
XFILLER_0_126_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13258_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[109\] _07610_ keymem.key_mem\[14\]\[109\]
+ _07666_ _08752_ sky130_fd_sc_hd__a22o_2
XFILLER_0_177_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_228 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12209_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[11\] _07683_ keymem.key_mem\[3\]\[11\]
+ _07603_ _07801_ sky130_fd_sc_hd__a22o_2
X_13189_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[102\] _07843_ keymem.key_mem\[2\]\[102\]
+ _07545_ _08690_ sky130_fd_sc_hd__a22o_2
XFILLER_0_97_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_209_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19805_ VGND VPWR VPWR VGND _05303_ keymem.key_mem\[11\]\[61\] _03162_ _05312_ sky130_fd_sc_hd__mux2_2
XFILLER_0_236_442 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17997_ VGND VPWR VGND VPWR _03929_ _03792_ _03795_ _03859_ _03727_ _03930_ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_97_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_58_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_236_486 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_172_2_Right_244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16948_ VGND VPWR VGND VPWR _03079_ _09513_ _10366_ key[53] sky130_fd_sc_hd__o21a_2
X_19736_ VGND VPWR VPWR VGND _05270_ keymem.key_mem\[11\]\[28\] _02787_ _05276_ sky130_fd_sc_hd__mux2_2
XFILLER_0_126_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16879_ VGND VPWR _00058_ _03016_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_223_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19667_ VGND VPWR _00625_ _05237_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_250_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18618_ VGND VPWR _04487_ _03957_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_232_692 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_172_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19598_ VGND VPWR VGND VPWR _05201_ keymem.key_mem_we _03435_ _05187_ _00592_ sky130_fd_sc_hd__a31o_2
XFILLER_0_19_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18549_ VGND VPWR _04425_ _03977_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_73_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1280 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_191_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21560_ VGND VPWR _01511_ _06244_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_34_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_929 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_56_970 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20511_ VGND VPWR VPWR VGND _05680_ _10661_ keymem.key_mem\[8\]\[8\] _05687_ sky130_fd_sc_hd__mux2_2
XFILLER_0_142_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21491_ VGND VPWR VPWR VGND _06196_ _03355_ keymem.key_mem\[5\]\[83\] _06208_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_834 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_439 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23230_ VGND VPWR _07118_ enc_block.block_w3_reg\[27\] enc_block.block_w0_reg\[19\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20442_ VGND VPWR VPWR VGND _05649_ _03518_ keymem.key_mem\[9\]\[104\] _05650_ sky130_fd_sc_hd__mux2_2
XFILLER_0_42_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_67_1173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23161_ VGND VPWR VGND VPWR _03582_ _02398_ _03584_ _07065_ sky130_fd_sc_hd__a21o_2
X_20373_ VGND VPWR _00955_ _05613_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_3_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_336 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_31_859 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_105_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22112_ VGND VPWR _01768_ _06539_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_144_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23092_ VGND VPWR VGND VPWR _02266_ _07021_ _07010_ keymem.prev_key1_reg\[89\] sky130_fd_sc_hd__o21a_2
XFILLER_0_3_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_282 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_80_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22043_ VGND VPWR VGND VPWR _06503_ keymem.key_mem_we _03356_ _06498_ _01735_ sky130_fd_sc_hd__a31o_2
XFILLER_0_45_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25802_ keymem.prev_key1_reg\[118\] clk _02295_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_23994_ VGND VPWR VPWR VGND clk _00487_ reset_n keymem.key_mem\[13\]\[115\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_138_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25733_ keymem.prev_key1_reg\[49\] clk _02226_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_214_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_202_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22945_ VGND VPWR VPWR VGND _02206_ _02798_ _02810_ _06925_ _06934_ sky130_fd_sc_hd__o31a_2
XFILLER_0_138_1167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_1117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_214_1022 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25664_ VGND VPWR VPWR VGND clk _02157_ reset_n keymem.key_mem\[0\]\[121\] sky130_fd_sc_hd__dfrtp_2
X_22876_ VGND VPWR _06891_ _06890_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_116_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_151_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24615_ VGND VPWR VPWR VGND clk _01108_ reset_n keymem.key_mem\[8\]\[96\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_112_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21827_ VGND VPWR _01637_ _06385_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_65_200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_91_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25595_ VGND VPWR VPWR VGND clk _02088_ reset_n keymem.key_mem\[0\]\[52\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_151_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_319 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_52_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_210_397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12560_ VGND VPWR VGND VPWR _08123_ _07737_ keymem.key_mem\[1\]\[40\] _08120_ _08122_
+ sky130_fd_sc_hd__a211o_2
X_24546_ VGND VPWR VPWR VGND clk _01039_ reset_n keymem.key_mem\[8\]\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_65_244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21758_ VGND VPWR _01604_ _06349_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_19_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20709_ VGND VPWR _01114_ _05790_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_80_214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12491_ VGND VPWR VGND VPWR _07691_ keymem.key_mem\[3\]\[34\] _08057_ _08059_ _08060_
+ _07663_ sky130_fd_sc_hd__a2111o_2
X_24477_ VGND VPWR VPWR VGND clk _00970_ reset_n keymem.key_mem\[9\]\[86\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_34_620 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21689_ VGND VPWR _01571_ _06313_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_34_631 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_266_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14230_ VGND VPWR VGND VPWR _09140_ _09033_ _09121_ _09701_ sky130_fd_sc_hd__a21o_2
XFILLER_0_46_491 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23428_ VGND VPWR _07296_ _04223_ _02327_ _07096_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_80_269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_199_Left_466 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_116_390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14161_ VPWR VGND VPWR VGND _09632_ keymem.prev_key1_reg\[65\] sky130_fd_sc_hd__inv_2
XFILLER_0_46_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23359_ _07233_ _07235_ _04103_ _07234_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_123_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13112_ VPWR VGND VPWR VGND _08620_ keymem.key_mem\[11\]\[94\] _08011_ keymem.key_mem\[8\]\[94\]
+ _08265_ _08621_ sky130_fd_sc_hd__a221o_2
XFILLER_0_127_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_131_360 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14092_ VGND VPWR _09563_ _09562_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_60_Left_328 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_131_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_123_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17920_ VGND VPWR VPWR VGND _03874_ _03877_ keymem.prev_key0_reg\[97\] _03878_ sky130_fd_sc_hd__mux2_2
X_13043_ VGND VPWR enc_block.round_key\[87\] _08558_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25029_ VGND VPWR VPWR VGND clk _01522_ reset_n keymem.key_mem\[5\]\[126\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_197_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17851_ VGND VPWR _00216_ _03830_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_219_987 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_203_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_272 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16802_ VGND VPWR _00051_ _02946_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17782_ VGND VPWR VPWR VGND _03719_ key[182] keymem.prev_key1_reg\[54\] _03783_ sky130_fd_sc_hd__mux2_2
X_14994_ VPWR VGND VPWR VGND _10457_ _10445_ _10444_ _10419_ _10458_ sky130_fd_sc_hd__or4_2
XFILLER_0_205_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19521_ VPWR VGND keymem.key_mem\[12\]\[56\] _05161_ _05158_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16733_ VGND VPWR _02884_ _09863_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13945_ VPWR VGND VPWR VGND _09261_ _09245_ _09266_ _09254_ _09417_ sky130_fd_sc_hd__or4_2
XFILLER_0_205_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19452_ VPWR VGND keymem.key_mem\[12\]\[24\] _05124_ _05116_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16664_ VGND VPWR VGND VPWR _02586_ _02572_ keymem.rcon_logic.tmp_rcon\[7\] _02818_
+ sky130_fd_sc_hd__a21o_2
X_13876_ VGND VPWR _09348_ _09347_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_134_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_202_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_198_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15615_ VPWR VGND VPWR VGND _11073_ _10504_ _10593_ sky130_fd_sc_hd__or2_2
X_18403_ VGND VPWR _04294_ _03981_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_243_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_70_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12827_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[66\] _07632_ keymem.key_mem\[1\]\[66\]
+ _07714_ _08364_ sky130_fd_sc_hd__a22o_2
X_19383_ VPWR VGND keymem.key_mem_we _05083_ _03647_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16595_ VGND VPWR _02752_ keymem.prev_key0_reg\[27\] _02751_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_232_1188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18334_ VPWR VGND VGND VPWR _04232_ _04233_ _04190_ sky130_fd_sc_hd__nor2_2
X_15546_ VPWR VGND VPWR VGND _10999_ _11004_ _11001_ _10637_ _11005_ sky130_fd_sc_hd__or4_2
XFILLER_0_70_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_31_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12758_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[59\] _07608_ keymem.key_mem\[11\]\[59\]
+ _07599_ _08302_ sky130_fd_sc_hd__a22o_2
XFILLER_0_267_1229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_210_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18265_ VPWR VGND VGND VPWR _04169_ _04170_ _04041_ sky130_fd_sc_hd__nor2_2
XFILLER_0_56_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11709_ VGND VPWR result[21] _07418_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15477_ VGND VPWR VGND VPWR _10644_ _10485_ _10595_ _10515_ _10475_ _10937_ sky130_fd_sc_hd__o32a_2
XFILLER_0_71_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12689_ VGND VPWR enc_block.round_key\[52\] _08239_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_210_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_115_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17216_ VGND VPWR VGND VPWR _03321_ _03152_ key[207] _03317_ _03320_ sky130_fd_sc_hd__a211o_2
X_14428_ VPWR VGND VPWR VGND _09897_ _09327_ _09582_ sky130_fd_sc_hd__or2_2
X_18196_ VPWR VGND VPWR VGND _04107_ _03970_ _02344_ sky130_fd_sc_hd__or2_2
XFILLER_0_126_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_804 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_245_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_24_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1313 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17147_ VPWR VGND VPWR VGND _03258_ _03257_ _03255_ _02497_ _03254_ _03259_ sky130_fd_sc_hd__a221o_2
X_14359_ VPWR VGND VGND VPWR _09050_ _09829_ _09138_ sky130_fd_sc_hd__nor2_2
XFILLER_0_40_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17078_ VGND VPWR keymem.prev_key0_reg\[65\] _09710_ _03197_ _09711_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_204_1224 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_180_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16029_ VPWR VGND VGND VPWR _11283_ _11484_ _11239_ sky130_fd_sc_hd__nor2_2
XFILLER_0_141_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1025 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_23_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_946 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_173_2_Right_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_97_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_776 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19719_ VGND VPWR VPWR VGND _05259_ keymem.key_mem\[11\]\[20\] _02480_ _05267_ sky130_fd_sc_hd__mux2_2
XFILLER_0_197_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20991_ VGND VPWR VPWR VGND _05934_ _05041_ keymem.key_mem\[7\]\[104\] _05943_ sky130_fd_sc_hd__mux2_2
XFILLER_0_211_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_215_1320 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_250_1211 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22730_ VGND VPWR VPWR VGND _06822_ keymem.key_mem\[0\]\[60\] _03150_ _06830_ sky130_fd_sc_hd__mux2_2
XFILLER_0_189_371 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_189_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_215_1364 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_212_Left_479 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22661_ VGND VPWR VPWR VGND _06798_ keymem.key_mem\[0\]\[19\] _02410_ _06802_ sky130_fd_sc_hd__mux2_2
XFILLER_0_220_695 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24400_ VGND VPWR VPWR VGND clk _00893_ reset_n keymem.key_mem\[9\]\[9\] sky130_fd_sc_hd__dfrtp_2
X_21612_ VPWR VGND VGND VPWR _06259_ _06273_ keymem.key_mem\[4\]\[11\] sky130_fd_sc_hd__nor2_2
X_25380_ VGND VPWR VPWR VGND clk _01873_ reset_n keymem.key_mem\[2\]\[93\] sky130_fd_sc_hd__dfrtp_2
X_22592_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[104\] _06775_ _06774_ _05041_ _02012_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_34_1194 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_8_842 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_266 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_104_1_Left_371 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_164_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24331_ VGND VPWR VPWR VGND clk _00824_ reset_n keymem.key_mem\[10\]\[68\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_1424 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21543_ VGND VPWR _01503_ _06235_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_28_491 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_105_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_209_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21474_ VGND VPWR _06199_ _03279_ _01470_ _06114_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_24262_ VGND VPWR VPWR VGND clk _00755_ reset_n keymem.key_mem\[11\]\[127\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_7_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_69_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23213_ _07101_ _07103_ _04064_ _07102_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_20425_ VGND VPWR VPWR VGND _05638_ _03466_ keymem.key_mem\[9\]\[96\] _05641_ sky130_fd_sc_hd__mux2_2
X_24193_ VGND VPWR VPWR VGND clk _00686_ reset_n keymem.key_mem\[11\]\[58\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_30_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_221_Left_488 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23144_ VGND VPWR _02284_ _07055_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20356_ VGND VPWR VPWR VGND _05602_ _03184_ keymem.key_mem\[9\]\[63\] _05605_ sky130_fd_sc_hd__mux2_2
XFILLER_0_259_353 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_109_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_248_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23075_ VGND VPWR VGND VPWR _02258_ _07012_ _07010_ keymem.prev_key1_reg\[81\] sky130_fd_sc_hd__o21a_2
XFILLER_0_41_1121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20287_ VGND VPWR _00914_ _05568_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_228_751 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22026_ VGND VPWR _06494_ _06402_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_216_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_196_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_76_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_243_776 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23977_ VGND VPWR VPWR VGND clk _00470_ reset_n keymem.key_mem\[13\]\[98\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_215_489 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11991_ VPWR VGND VGND VPWR _07548_ _07594_ _07554_ sky130_fd_sc_hd__nor2_2
X_13730_ _09184_ _09202_ _09039_ _09046_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_230_Left_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25716_ keymem.prev_key1_reg\[32\] clk _02209_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22928_ VGND VPWR VGND VPWR _06923_ _02676_ _06891_ _02687_ _06892_ sky130_fd_sc_hd__a211o_2
XFILLER_0_85_306 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13661_ VGND VPWR VPWR VGND _09058_ _09017_ _08958_ _09133_ sky130_fd_sc_hd__or3_2
XFILLER_0_97_188 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25647_ VGND VPWR VPWR VGND clk _02140_ reset_n keymem.key_mem\[0\]\[104\] sky130_fd_sc_hd__dfrtp_2
X_22859_ VGND VPWR _06878_ _06877_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15400_ VGND VPWR VGND VPWR _10850_ _10860_ _10861_ _10844_ _10855_ sky130_fd_sc_hd__nor4_2
XFILLER_0_13_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12612_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[45\] _07771_ keymem.key_mem\[9\]\[45\]
+ _07592_ _08170_ sky130_fd_sc_hd__a22o_2
XFILLER_0_155_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16380_ VPWR VGND VPWR VGND _02541_ _02543_ _02539_ _02540_ sky130_fd_sc_hd__or3b_2
X_13592_ VGND VPWR VGND VPWR _09064_ _09026_ _09025_ keymem.prev_key1_reg\[0\] _08956_
+ _08943_ sky130_fd_sc_hd__a32o_2
X_25578_ VGND VPWR VPWR VGND clk _02071_ reset_n keymem.key_mem\[0\]\[35\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15331_ VPWR VGND VPWR VGND _10715_ _10792_ _10789_ _10643_ _10793_ sky130_fd_sc_hd__or4_2
XFILLER_0_38_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12543_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[39\] _07918_ keymem.key_mem\[4\]\[39\]
+ _07913_ _08107_ sky130_fd_sc_hd__a22o_2
X_24529_ VGND VPWR VPWR VGND clk _01022_ reset_n keymem.key_mem\[8\]\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26_439 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_87_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18050_ VPWR VGND VGND VPWR _07374_ _03972_ _08923_ sky130_fd_sc_hd__nor2_2
X_15262_ VGND VPWR VGND VPWR _10588_ _10547_ _10519_ _10725_ sky130_fd_sc_hd__a21o_2
X_12474_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[32\] _07536_ _08044_ _08040_ _08045_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_87_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17001_ VPWR VGND VPWR VGND _03127_ key[186] _10322_ sky130_fd_sc_hd__or2_2
X_14213_ VGND VPWR _09684_ _09683_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15193_ VPWR VGND VGND VPWR _09796_ _10657_ key[8] sky130_fd_sc_hd__nor2_2
XFILLER_0_22_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14144_ VGND VPWR VGND VPWR _09614_ _09613_ _09615_ _09612_ _09611_ sky130_fd_sc_hd__nand4_2
XFILLER_0_123_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18952_ VGND VPWR _04788_ _03949_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14075_ VPWR VGND VPWR VGND _09546_ _09545_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13026_ VPWR VGND VPWR VGND _08542_ keymem.key_mem\[14\]\[86\] _08003_ keymem.key_mem\[8\]\[86\]
+ _07655_ _08543_ sky130_fd_sc_hd__a221o_2
X_17903_ VPWR VGND VPWR VGND _03866_ _03865_ keymem.prev_key0_reg\[91\] _03788_ _00232_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_20_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18883_ VGND VPWR VPWR VGND _04600_ enc_block.block_w2_reg\[13\] _04125_ _04726_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_158_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_148_2_Left_619 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17834_ VGND VPWR VGND VPWR _03243_ keymem.prev_key1_reg\[70\] _03819_ _03818_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_98_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_26 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14977_ VGND VPWR VPWR VGND _10440_ _10409_ _10439_ _10441_ sky130_fd_sc_hd__or3_2
X_17765_ VGND VPWR _00187_ _03773_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19504_ VGND VPWR VPWR VGND _05151_ _04950_ keymem.key_mem\[12\]\[48\] _05152_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13928_ VPWR VGND VPWR VGND _09280_ _09309_ _09321_ _09338_ _09400_ sky130_fd_sc_hd__or4_2
X_16716_ VGND VPWR VPWR VGND _02867_ _02868_ _08931_ _02342_ _09508_ sky130_fd_sc_hd__a31oi_2
X_17696_ VGND VPWR _03727_ _03672_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_16_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19435_ VGND VPWR VGND VPWR _05114_ keymem.key_mem_we _11447_ _05109_ _00516_ sky130_fd_sc_hd__a31o_2
X_16647_ VGND VPWR keymem.prev_key1_reg\[125\] _02799_ _02802_ _02800_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_13859_ VGND VPWR _09331_ _09299_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_76_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_31_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_639 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19366_ VGND VPWR VPWR VGND _05067_ _05071_ keymem.key_mem\[13\]\[118\] _05072_ sky130_fd_sc_hd__mux2_2
X_16578_ VGND VPWR keymem.prev_key1_reg\[90\] _02733_ _02736_ _02734_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_32_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_267_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15529_ VPWR VGND VGND VPWR _10467_ _10545_ _10988_ _10481_ _10534_ sky130_fd_sc_hd__o22ai_2
X_18317_ VPWR VGND VPWR VGND _04217_ enc_block.block_w2_reg\[13\] enc_block.block_w2_reg\[14\]
+ sky130_fd_sc_hd__or2_2
XFILLER_0_123_76 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_169_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19297_ VGND VPWR _05025_ _04876_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_32_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18248_ VPWR VGND VGND VPWR _04154_ _04079_ _04153_ sky130_fd_sc_hd__nand2_2
XFILLER_0_66_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18179_ VGND VPWR _04091_ _04088_ _04090_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_167_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_1121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20210_ VGND VPWR VPWR VGND _05388_ _03647_ keymem.key_mem\[10\]\[124\] _05526_ sky130_fd_sc_hd__mux2_2
X_21190_ VGND VPWR VPWR VGND _06040_ _03234_ keymem.key_mem\[6\]\[69\] _06049_ sky130_fd_sc_hd__mux2_2
XFILLER_0_141_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_312 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_145_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20141_ VGND VPWR VPWR VGND _05482_ _03427_ keymem.key_mem\[10\]\[91\] _05490_ sky130_fd_sc_hd__mux2_2
XFILLER_0_0_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20072_ VGND VPWR VPWR VGND _05446_ _03130_ keymem.key_mem\[10\]\[58\] _05454_ sky130_fd_sc_hd__mux2_2
XFILLER_0_42_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23900_ VGND VPWR VPWR VGND clk _00393_ reset_n keymem.key_mem\[13\]\[21\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24880_ VGND VPWR VPWR VGND clk _01373_ reset_n keymem.key_mem\[6\]\[105\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_256_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_905 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23831_ VGND VPWR VPWR VGND clk _00324_ reset_n enc_block.block_w1_reg\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_174_2_Right_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_1201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23762_ keymem.prev_key0_reg\[118\] clk _00259_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_79_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20974_ VGND VPWR _05934_ _05819_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_73_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25501_ VGND VPWR VPWR VGND clk _01994_ reset_n keymem.key_mem\[1\]\[86\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_67_317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22713_ VGND VPWR _06822_ _06778_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_117_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23693_ keymem.prev_key0_reg\[49\] clk _00190_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_113_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1074 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_220_481 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25432_ VGND VPWR VPWR VGND clk _01925_ reset_n keymem.key_mem\[1\]\[17\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_194_2_Left_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_53_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22644_ VGND VPWR _02046_ _06793_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_187_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_333 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_63_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_113_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_203 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_737 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25363_ VGND VPWR VPWR VGND clk _01856_ reset_n keymem.key_mem\[2\]\[76\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_187_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22575_ VGND VPWR VPWR VGND _06701_ keymem.key_mem\[1\]\[92\] _03435_ _06771_ sky130_fd_sc_hd__mux2_2
XFILLER_0_8_661 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24314_ VGND VPWR VPWR VGND clk _00807_ reset_n keymem.key_mem\[10\]\[51\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_263_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21526_ VGND VPWR _01495_ _06226_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_228_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25294_ VGND VPWR VPWR VGND clk _01787_ reset_n keymem.key_mem\[2\]\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_263_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24245_ VGND VPWR VPWR VGND clk _00738_ reset_n keymem.key_mem\[11\]\[110\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_160_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21457_ VGND VPWR _01462_ _06190_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_224_1419 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_259_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_802 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20408_ VGND VPWR VPWR VGND _05627_ _03401_ keymem.key_mem\[9\]\[88\] _05632_ sky130_fd_sc_hd__mux2_2
X_12190_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[10\] _07782_ keymem.key_mem\[11\]\[10\]
+ _07781_ _07783_ sky130_fd_sc_hd__a22o_2
X_24176_ VGND VPWR VPWR VGND clk _00669_ reset_n keymem.key_mem\[11\]\[41\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_266_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21388_ VGND VPWR _01429_ _06154_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_124_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23127_ VGND VPWR VPWR VGND _07032_ _07043_ keymem.prev_key1_reg\[102\] _07044_ sky130_fd_sc_hd__mux2_2
X_20339_ VGND VPWR VPWR VGND _05591_ _03099_ keymem.key_mem\[9\]\[55\] _05596_ sky130_fd_sc_hd__mux2_2
XFILLER_0_124_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23058_ VGND VPWR VGND VPWR _07001_ _03794_ _03285_ _07002_ sky130_fd_sc_hd__a21o_2
XFILLER_0_21_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14900_ VPWR VGND VPWR VGND _10330_ _10364_ _10363_ _09516_ _10365_ sky130_fd_sc_hd__or4_2
X_22009_ VGND VPWR VGND VPWR _06485_ keymem.key_mem_we _03217_ _06475_ _01719_ sky130_fd_sc_hd__a31o_2
X_15880_ VGND VPWR _11336_ _11262_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14831_ VPWR VGND VPWR VGND _10123_ _10295_ _10296_ _09877_ _10294_ sky130_fd_sc_hd__or4b_2
XFILLER_0_235_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_426 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17550_ VGND VPWR _00131_ _03614_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14762_ VPWR VGND VPWR VGND _09692_ _10227_ _09947_ _09093_ _10228_ sky130_fd_sc_hd__or4_2
XFILLER_0_231_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11974_ VGND VPWR _07577_ _07576_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_230_256 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16501_ VGND VPWR _02662_ _09863_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_212_960 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13713_ VGND VPWR _09185_ _09041_ _09039_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_17481_ VPWR VGND VPWR VGND _03554_ _09534_ _03552_ key[238] _03527_ _03555_ sky130_fd_sc_hd__a221o_2
X_14693_ VPWR VGND VPWR VGND _10159_ _10160_ _09675_ _10158_ sky130_fd_sc_hd__or3b_2
XFILLER_0_224_64 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16432_ VGND VPWR VGND VPWR _02592_ _02591_ _02594_ _02593_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_131_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19220_ VGND VPWR VPWR VGND _04951_ _04977_ keymem.key_mem\[13\]\[66\] _04978_ sky130_fd_sc_hd__mux2_2
X_13644_ VGND VPWR _09116_ _09115_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_85_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_128_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19151_ VPWR VGND keymem.key_mem_we _04935_ _02955_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_2_1029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16363_ VPWR VGND VPWR VGND _02519_ _02525_ _02523_ _02434_ _02526_ sky130_fd_sc_hd__or4_2
X_13575_ VPWR VGND VGND VPWR _09010_ _09047_ _08958_ sky130_fd_sc_hd__nor2_2
XFILLER_0_211_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_236 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_759 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18102_ VPWR VGND VPWR VGND _04020_ _03992_ _04018_ enc_block.block_w0_reg\[3\] _03976_
+ _00277_ sky130_fd_sc_hd__a221o_2
XFILLER_0_26_247 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15314_ VGND VPWR VGND VPWR _10674_ _10776_ _10572_ _10569_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_240_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12526_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[37\] _07565_ keymem.key_mem\[1\]\[37\]
+ _07855_ _08092_ sky130_fd_sc_hd__a22o_2
X_19082_ VGND VPWR VPWR VGND _04877_ _04894_ keymem.key_mem\[13\]\[11\] _04895_ sky130_fd_sc_hd__mux2_2
X_16294_ VPWR VGND VGND VPWR _02435_ _02443_ _02457_ _02458_ sky130_fd_sc_hd__nor3_2
XFILLER_0_136_282 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18033_ VGND VPWR VPWR VGND enc_block.sword_ctr_inc enc_block.enc_ctrl_reg\[3\] _03955_
+ _07374_ _07381_ sky130_fd_sc_hd__o211a_2
XFILLER_0_240_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15245_ VPWR VGND VGND VPWR _10498_ _10504_ _10708_ _10635_ _10588_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_48_1149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12457_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[31\] _07586_ keymem.key_mem\[1\]\[31\]
+ _07624_ _08029_ sky130_fd_sc_hd__a22o_2
XFILLER_0_169_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15176_ VPWR VGND VGND VPWR _10639_ _10640_ _10565_ sky130_fd_sc_hd__nor2_2
XFILLER_0_111_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12388_ VPWR VGND VPWR VGND _07965_ keymem.key_mem\[5\]\[25\] _07811_ keymem.key_mem\[13\]\[25\]
+ _07622_ _07966_ sky130_fd_sc_hd__a221o_2
XFILLER_0_1_347 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14127_ VPWR VGND VPWR VGND _09591_ _09597_ _09592_ _09590_ _09598_ sky130_fd_sc_hd__or4_2
XFILLER_0_50_795 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19984_ VGND VPWR VPWR VGND _05400_ _11447_ keymem.key_mem\[10\]\[16\] _05408_ sky130_fd_sc_hd__mux2_2
X_18935_ VPWR VGND _04772_ enc_block.block_w0_reg\[10\] enc_block.block_w1_reg\[3\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_14058_ VGND VPWR VPWR VGND _09511_ _09530_ _09528_ _09526_ _09527_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_185_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_197_1153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13009_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[84\] _07578_ keymem.key_mem\[8\]\[84\]
+ _07903_ _08528_ sky130_fd_sc_hd__a22o_2
XFILLER_0_182_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18866_ VPWR VGND _04710_ _04635_ enc_block.block_w1_reg\[4\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_98_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17817_ VGND VPWR VPWR VGND _03777_ _03806_ keymem.prev_key0_reg\[65\] _03807_ sky130_fd_sc_hd__mux2_2
XFILLER_0_206_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18797_ VGND VPWR _04648_ enc_block.block_w1_reg\[4\] _04647_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_265_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17748_ VGND VPWR _03763_ _03674_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_171_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17679_ VGND VPWR VPWR VGND _03703_ _03715_ keymem.prev_key0_reg\[18\] _03716_ sky130_fd_sc_hd__mux2_2
XFILLER_0_134_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_174_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_251_1394 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19418_ VGND VPWR VGND VPWR _05105_ keymem.key_mem_we _10662_ _05093_ _00508_ sky130_fd_sc_hd__a31o_2
X_20690_ VGND VPWR _01105_ _05780_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_64_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19349_ VPWR VGND keymem.key_mem_we _05060_ _03573_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_17_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1255 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_150_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22360_ VGND VPWR VPWR VGND _06669_ _03525_ keymem.key_mem\[2\]\[105\] _06671_ sky130_fd_sc_hd__mux2_2
XFILLER_0_26_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21311_ VGND VPWR VPWR VGND _05971_ _03668_ keymem.key_mem\[6\]\[127\] _06112_ sky130_fd_sc_hd__mux2_2
XFILLER_0_87_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22291_ VGND VPWR VPWR VGND _06634_ _03259_ keymem.key_mem\[2\]\[72\] _06635_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_32_239 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_142_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21242_ VGND VPWR _06076_ _05970_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24030_ VGND VPWR VPWR VGND clk _00523_ reset_n keymem.key_mem\[12\]\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_206_1138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_762 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_206_1149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_29_1060 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_182_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21173_ VGND VPWR _06040_ _05970_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_159_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_106_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20124_ VGND VPWR VPWR VGND _05469_ _03356_ keymem.key_mem\[10\]\[83\] _05481_ sky130_fd_sc_hd__mux2_2
XFILLER_0_141_1174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_256_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20055_ VGND VPWR VPWR VGND _05435_ _03056_ keymem.key_mem\[10\]\[50\] _05445_ sky130_fd_sc_hd__mux2_2
X_24932_ VGND VPWR VPWR VGND clk _01425_ reset_n keymem.key_mem\[5\]\[29\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24863_ VGND VPWR VPWR VGND clk _01356_ reset_n keymem.key_mem\[6\]\[88\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23814_ VGND VPWR VPWR VGND clk _00307_ reset_n enc_block.sword_ctr_reg\[1\] sky130_fd_sc_hd__dfrtp_2
X_24794_ VGND VPWR VPWR VGND clk _01287_ reset_n keymem.key_mem\[6\]\[19\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_175_2_Right_247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_217_1278 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_201_919 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23745_ keymem.prev_key0_reg\[101\] clk _00242_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_67_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20957_ VGND VPWR VGND VPWR _05925_ keymem.key_mem_we _03393_ _05916_ _01227_ sky130_fd_sc_hd__a31o_2
XFILLER_0_191_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11690_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[12\] dec_new_block\[12\]
+ _07409_ sky130_fd_sc_hd__mux2_2
XFILLER_0_67_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23676_ keymem.prev_key0_reg\[32\] clk _00173_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20888_ VGND VPWR VPWR VGND _05880_ _04963_ keymem.key_mem\[7\]\[55\] _05889_ sky130_fd_sc_hd__mux2_2
X_25415_ VGND VPWR VPWR VGND clk _01908_ reset_n keymem.key_mem\[1\]\[0\] sky130_fd_sc_hd__dfrtp_2
X_22627_ VGND VPWR _02039_ _06783_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25346_ VGND VPWR VPWR VGND clk _01839_ reset_n keymem.key_mem\[2\]\[59\] sky130_fd_sc_hd__dfrtp_2
X_13360_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[119\] _07666_ keymem.key_mem\[4\]\[119\]
+ _08077_ _08844_ sky130_fd_sc_hd__a22o_2
XFILLER_0_180_325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_88_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22558_ VGND VPWR VPWR VGND _06750_ keymem.key_mem\[1\]\[82\] _03347_ _06764_ sky130_fd_sc_hd__mux2_2
XFILLER_0_148_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12311_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[19\] _07818_ keymem.key_mem\[12\]\[19\]
+ _07894_ _07895_ sky130_fd_sc_hd__a22o_2
X_21509_ VGND VPWR _01487_ _06217_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_23_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25277_ VGND VPWR VPWR VGND clk _01770_ reset_n keymem.key_mem\[3\]\[118\] sky130_fd_sc_hd__dfrtp_2
X_13291_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[112\] _07742_ keymem.key_mem\[12\]\[112\]
+ _07787_ _08782_ sky130_fd_sc_hd__a22o_2
XFILLER_0_49_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22489_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[41\] _06707_ _06706_ _04937_ _01949_
+ sky130_fd_sc_hd__a22o_2
X_15030_ VPWR VGND VPWR VGND _10424_ _10445_ _10430_ _10443_ _10494_ sky130_fd_sc_hd__or4_2
X_24228_ VGND VPWR VPWR VGND clk _00721_ reset_n keymem.key_mem\[11\]\[93\] sky130_fd_sc_hd__dfrtp_2
X_12242_ VGND VPWR enc_block.round_key\[13\] _07831_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_239_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24159_ VGND VPWR VPWR VGND clk _00652_ reset_n keymem.key_mem\[11\]\[24\] sky130_fd_sc_hd__dfrtp_2
X_12173_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[9\] _07595_ keymem.key_mem\[9\]\[9\]
+ _07591_ _07767_ sky130_fd_sc_hd__a22o_2
XFILLER_0_48_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_816 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_182 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_257_1003 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16981_ VGND VPWR _03109_ _03108_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_219_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18720_ VPWR VGND VGND VPWR _04578_ _04434_ _04577_ sky130_fd_sc_hd__nand2_2
XFILLER_0_263_646 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_235_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_159_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15932_ VGND VPWR VGND VPWR _11388_ _11386_ _11253_ _11311_ _11205_ _11387_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_95_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15863_ VPWR VGND VPWR VGND _11265_ _11221_ _11179_ _11166_ _11319_ sky130_fd_sc_hd__or4_2
X_18651_ VGND VPWR _04517_ _04515_ _04516_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_239_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14814_ VGND VPWR VGND VPWR _10280_ _10277_ _10272_ _10092_ _10279_ sky130_fd_sc_hd__o211ai_2
X_17602_ VPWR VGND VGND VPWR keylen _03658_ _03659_ _03660_ sky130_fd_sc_hd__nor3_2
XFILLER_0_204_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_157_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15794_ VGND VPWR _11250_ _11249_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18582_ VPWR VGND VPWR VGND _04455_ _04307_ _04453_ sky130_fd_sc_hd__or2_2
XFILLER_0_58_103 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14745_ VPWR VGND VPWR VGND _09994_ _10210_ _10211_ _09846_ _09963_ sky130_fd_sc_hd__or4b_2
X_17533_ VGND VPWR VGND VPWR _03152_ key[245] _03599_ _03600_ sky130_fd_sc_hd__a21o_2
XFILLER_0_54_1142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11957_ VGND VPWR _07560_ _07559_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_59_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1186 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17464_ VGND VPWR VPWR VGND _03029_ _10963_ key[108] _03540_ sky130_fd_sc_hd__mux2_2
XFILLER_0_46_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1028 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14676_ VPWR VGND _10143_ _10142_ keymem.prev_key1_reg\[69\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_11888_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[15\] dec_new_block\[111\]
+ _07508_ sky130_fd_sc_hd__mux2_2
XFILLER_0_39_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16415_ VGND VPWR VGND VPWR _11370_ _11318_ _02577_ _11298_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_7_907 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_251_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19203_ VGND VPWR _04968_ _04877_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13627_ VGND VPWR _09099_ _09098_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17395_ VGND VPWR VPWR VGND _03467_ keymem.key_mem\[14\]\[98\] _03480_ _03481_ sky130_fd_sc_hd__mux2_2
XFILLER_0_156_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_854 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_55_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16346_ VPWR VGND VPWR VGND _02507_ _02508_ _02509_ _11488_ _11562_ sky130_fd_sc_hd__or4b_2
XFILLER_0_67_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19134_ VGND VPWR _04924_ _04877_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13558_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[3\] _08956_ _09030_ _08943_ _08961_
+ _08962_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_15_729 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_246_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12509_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[36\] _07838_ keymem.key_mem\[2\]\[36\]
+ _07816_ _08076_ sky130_fd_sc_hd__a22o_2
X_19065_ VPWR VGND keymem.key_mem\[13\]\[4\] _04885_ _04880_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16277_ VPWR VGND VGND VPWR _11307_ _11334_ _02441_ _11303_ _11385_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_28_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13489_ VPWR VGND VPWR VGND _08960_ _08948_ _08959_ _08945_ enc_block.block_w2_reg\[3\]
+ _08961_ sky130_fd_sc_hd__a221o_2
XFILLER_0_246_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15228_ VGND VPWR VGND VPWR _10527_ _10608_ _10691_ _10595_ sky130_fd_sc_hd__a21oi_2
X_18016_ VPWR VGND VGND VPWR _03942_ _00269_ _03941_ sky130_fd_sc_hd__nor2_2
XFILLER_0_23_762 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_2_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_924 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15159_ VGND VPWR VPWR VGND _10453_ _10477_ _10439_ _10623_ sky130_fd_sc_hd__or3_2
XFILLER_0_61_1124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_125_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_164 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_201_1035 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19967_ VGND VPWR _00764_ _05398_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18918_ VGND VPWR _04757_ _04754_ _04756_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_226_348 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_177_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19898_ VGND VPWR _00733_ _05360_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_113_1_Left_380 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_138_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18849_ _04693_ _04695_ _04692_ _04694_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_253_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1053 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_74_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_145_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_96_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21860_ VGND VPWR _06404_ _06403_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_214_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20811_ VGND VPWR VGND VPWR _05847_ keymem.key_mem_we _02410_ _05838_ _01159_ sky130_fd_sc_hd__a31o_2
X_21791_ VGND VPWR VPWR VGND _06366_ _03466_ keymem.key_mem\[4\]\[96\] _06367_ sky130_fd_sc_hd__mux2_2
XFILLER_0_72_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23530_ VGND VPWR VPWR VGND clk _00031_ reset_n keymem.key_mem\[14\]\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_158 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20742_ VGND VPWR VPWR VGND _05805_ _03607_ keymem.key_mem\[8\]\[118\] _05808_ sky130_fd_sc_hd__mux2_2
XFILLER_0_114_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_58_692 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23461_ VGND VPWR VGND VPWR _07325_ _04149_ _07093_ _07326_ enc_block.block_w3_reg\[26\]
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_174_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20673_ VGND VPWR _01097_ _05771_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25200_ VGND VPWR VPWR VGND clk _01693_ reset_n keymem.key_mem\[3\]\[41\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22412_ VGND VPWR _01909_ _06698_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23392_ VPWR VGND _07264_ enc_block.block_w1_reg\[10\] enc_block.block_w2_reg\[3\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_18_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_264_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25131_ VGND VPWR VPWR VGND clk _01624_ reset_n keymem.key_mem\[4\]\[100\] sky130_fd_sc_hd__dfrtp_2
X_22343_ VGND VPWR VPWR VGND _06658_ _03474_ keymem.key_mem\[2\]\[97\] _06662_ sky130_fd_sc_hd__mux2_2
XFILLER_0_225_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25062_ VGND VPWR VPWR VGND clk _01555_ reset_n keymem.key_mem\[4\]\[31\] sky130_fd_sc_hd__dfrtp_2
X_22274_ VGND VPWR VPWR VGND _06622_ _03193_ keymem.key_mem\[2\]\[64\] _06626_ sky130_fd_sc_hd__mux2_2
XFILLER_0_60_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24013_ VGND VPWR VPWR VGND clk _00506_ reset_n keymem.key_mem\[12\]\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_143_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21225_ VGND VPWR _01353_ _06067_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_130_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21156_ VGND VPWR _01320_ _06031_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_160_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_256_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20107_ VGND VPWR _05472_ _03279_ _00830_ _05402_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_217_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21087_ VGND VPWR VPWR VGND _05983_ _02479_ keymem.key_mem\[6\]\[20\] _05995_ sky130_fd_sc_hd__mux2_2
X_20038_ VGND VPWR _00797_ _05436_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_244_167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24915_ VGND VPWR VPWR VGND clk _01408_ reset_n keymem.key_mem\[5\]\[12\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_244_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24846_ VGND VPWR VPWR VGND clk _01339_ reset_n keymem.key_mem\[6\]\[71\] sky130_fd_sc_hd__dfrtp_2
X_12860_ VGND VPWR VGND VPWR _08394_ _07968_ keymem.key_mem\[9\]\[69\] _08390_ _08393_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_9_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11811_ VGND VPWR result[72] _07469_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_90_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_150_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12791_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[62\] _07645_ _08331_ _08325_ _08332_
+ sky130_fd_sc_hd__o22a_2
XPHY_EDGE_ROW_176_2_Right_248 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24777_ VGND VPWR VPWR VGND clk _01270_ reset_n keymem.key_mem\[6\]\[2\] sky130_fd_sc_hd__dfrtp_2
X_21989_ VGND VPWR VGND VPWR _06474_ keymem.key_mem_we _03130_ _06446_ _01710_ sky130_fd_sc_hd__a31o_2
XFILLER_0_154_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14530_ VPWR VGND VGND VPWR _09658_ _09222_ _09998_ _09160_ _09080_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_189_1417 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11742_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[6\] dec_new_block\[38\]
+ _07435_ sky130_fd_sc_hd__mux2_2
X_23728_ keymem.prev_key0_reg\[84\] clk _00225_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_90_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14461_ VGND VPWR _09930_ _09795_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_95_297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23659_ keymem.prev_key0_reg\[15\] clk _00156_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_11673_ VGND VPWR result[3] _07400_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_138_377 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16200_ _11291_ _02365_ _11338_ _11390_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_36_342 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13412_ VPWR VGND VPWR VGND _08890_ keymem.key_mem\[13\]\[124\] _07695_ keymem.key_mem\[1\]\[124\]
+ _07901_ _08891_ sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_189_1_Left_456 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17180_ VGND VPWR _03288_ _09541_ _00087_ _03287_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_70_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14392_ VGND VPWR _09862_ _09861_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_64_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_157_2_Left_628 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_153_358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16131_ VGND VPWR VGND VPWR _11311_ _11345_ _11375_ _11420_ _11585_ sky130_fd_sc_hd__o22a_2
X_25329_ VGND VPWR VPWR VGND clk _01822_ reset_n keymem.key_mem\[2\]\[42\] sky130_fd_sc_hd__dfrtp_2
X_13343_ VGND VPWR VGND VPWR _08829_ _07737_ keymem.key_mem\[1\]\[117\] _08826_ _08828_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_180_166 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_84_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16062_ VGND VPWR VGND VPWR _11284_ _11298_ _11278_ _11516_ _11412_ _11517_ sky130_fd_sc_hd__o32a_2
XFILLER_0_51_367 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_161_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13274_ VPWR VGND VPWR VGND _08766_ keymem.key_mem\[5\]\[110\] _07780_ keymem.key_mem\[14\]\[110\]
+ _07584_ _08767_ sky130_fd_sc_hd__a221o_2
XFILLER_0_59_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15013_ VGND VPWR _10477_ _10466_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_161_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12225_ VGND VPWR _07816_ _07732_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_62_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19821_ VGND VPWR _05320_ _03227_ _00696_ _05243_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_12156_ VGND VPWR enc_block.round_key\[7\] _07751_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_75_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19752_ VGND VPWR _00663_ _05284_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16964_ VGND VPWR VGND VPWR _02644_ _02643_ _10386_ _03093_ sky130_fd_sc_hd__a21o_2
XFILLER_0_224_808 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12087_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[4\] _07556_ keymem.key_mem\[2\]\[4\]
+ _07544_ _07686_ sky130_fd_sc_hd__a22o_2
X_18703_ VPWR VGND VGND VPWR _04563_ _04353_ _04562_ sky130_fd_sc_hd__nand2_2
XFILLER_0_263_476 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_194_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15915_ VPWR VGND VGND VPWR _11370_ _11371_ _11305_ sky130_fd_sc_hd__nor2_2
XFILLER_0_223_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19683_ VGND VPWR _00630_ _05248_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16895_ VGND VPWR VPWR VGND _03030_ _03031_ _09930_ _11160_ _11441_ sky130_fd_sc_hd__a31oi_2
X_18634_ VPWR VGND _04502_ _04501_ enc_block.round_key\[84\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_232_852 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15846_ VPWR VGND VPWR VGND _11192_ _11208_ _11197_ _11288_ _11302_ sky130_fd_sc_hd__or4_2
XFILLER_0_91_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_95_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_565 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_172_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_231_362 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_59_423 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18565_ VPWR VGND VPWR VGND _04439_ block[77] _04351_ enc_block.block_w3_reg\[13\]
+ _03954_ _04440_ sky130_fd_sc_hd__a221o_2
X_15777_ VGND VPWR _11233_ _11232_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12989_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[82\] _07673_ keymem.key_mem\[4\]\[82\]
+ _07692_ _08510_ sky130_fd_sc_hd__a22o_2
XFILLER_0_115_44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_172_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17516_ VPWR VGND VPWR VGND _03584_ _03582_ _02398_ key[243] _03527_ _03585_ sky130_fd_sc_hd__a221o_2
XFILLER_0_145_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14728_ VGND VPWR VPWR VGND _09864_ keymem.key_mem\[14\]\[5\] _10194_ _10195_ sky130_fd_sc_hd__mux2_2
X_18496_ VPWR VGND VPWR VGND _04377_ block[70] _04330_ enc_block.block_w0_reg\[6\]
+ _04276_ _04378_ sky130_fd_sc_hd__a221o_2
XFILLER_0_129_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14659_ VPWR VGND VGND VPWR _10126_ _10124_ _10125_ sky130_fd_sc_hd__nand2_2
X_17447_ VGND VPWR VPWR VGND _03467_ keymem.key_mem\[14\]\[105\] _03525_ _03526_ sky130_fd_sc_hd__mux2_2
XFILLER_0_27_364 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17378_ VPWR VGND VPWR VGND _03465_ _10902_ _03462_ key[224] _03366_ _03466_ sky130_fd_sc_hd__a221o_2
XFILLER_0_40_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_824 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_67_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19117_ VPWR VGND keymem.key_mem\[13\]\[27\] _04914_ _04903_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16329_ VGND VPWR VGND VPWR _02487_ _02486_ _02492_ keymem.prev_key1_reg\[85\] sky130_fd_sc_hd__a21oi_2
XFILLER_0_28_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_2_Right_210 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19048_ VGND VPWR _04873_ enc_block.round_key\[63\] _04872_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_242_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1030 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_242_1168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21010_ VGND VPWR VPWR VGND _05945_ _05060_ keymem.key_mem\[7\]\[113\] _05953_ sky130_fd_sc_hd__mux2_2
XFILLER_0_10_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_227_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_227_646 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_199_1089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_220_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22961_ VGND VPWR VGND VPWR _02907_ _06891_ _06944_ _02912_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24700_ VGND VPWR VPWR VGND clk _01193_ reset_n keymem.key_mem\[7\]\[53\] sky130_fd_sc_hd__dfrtp_2
X_21912_ VGND VPWR VGND VPWR _06433_ keymem.key_mem_we _02608_ _06432_ _01674_ sky130_fd_sc_hd__a31o_2
XFILLER_0_65_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25680_ VGND VPWR VPWR VGND clk _02173_ reset_n keymem.round_ctr_reg\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22892_ VGND VPWR VGND VPWR _10826_ _10825_ _10834_ _06901_ sky130_fd_sc_hd__a21o_2
XFILLER_0_190_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24631_ VGND VPWR VPWR VGND clk _01124_ reset_n keymem.key_mem\[8\]\[112\] sky130_fd_sc_hd__dfrtp_2
X_21843_ VGND VPWR VPWR VGND _06388_ _03627_ keymem.key_mem\[4\]\[121\] _06394_ sky130_fd_sc_hd__mux2_2
XFILLER_0_179_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_151_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24562_ VGND VPWR VPWR VGND clk _01055_ reset_n keymem.key_mem\[8\]\[43\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_172_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21774_ VGND VPWR VPWR VGND _06355_ _03401_ keymem.key_mem\[4\]\[88\] _06358_ sky130_fd_sc_hd__mux2_2
XFILLER_0_19_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23513_ VGND VPWR VPWR VGND clk _00014_ reset_n keymem.key_mem\[14\]\[2\] sky130_fd_sc_hd__dfrtp_2
X_20725_ VGND VPWR VPWR VGND _05794_ _03555_ keymem.key_mem\[8\]\[110\] _05799_ sky130_fd_sc_hd__mux2_2
X_24493_ VGND VPWR VPWR VGND clk _00986_ reset_n keymem.key_mem\[9\]\[102\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_1078 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_135_325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23444_ VPWR VGND VGND VPWR _07192_ _07311_ _04240_ sky130_fd_sc_hd__nor2_2
XFILLER_0_149_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20656_ VGND VPWR VPWR VGND _05761_ _03306_ keymem.key_mem\[8\]\[77\] _05763_ sky130_fd_sc_hd__mux2_2
XFILLER_0_162_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_18_397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23375_ VGND VPWR _07249_ _07176_ _07248_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_162_166 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20587_ VGND VPWR VPWR VGND _05725_ _02998_ keymem.key_mem\[8\]\[44\] _05727_ sky130_fd_sc_hd__mux2_2
X_25114_ VGND VPWR VPWR VGND clk _01607_ reset_n keymem.key_mem\[4\]\[83\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_367 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22326_ VGND VPWR VPWR VGND _06647_ _03409_ keymem.key_mem\[2\]\[89\] _06653_ sky130_fd_sc_hd__mux2_2
XFILLER_0_21_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_225_1355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_60_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25045_ VGND VPWR VPWR VGND clk _01538_ reset_n keymem.key_mem\[4\]\[14\] sky130_fd_sc_hd__dfrtp_2
X_22257_ VGND VPWR VPWR VGND _06611_ _03108_ keymem.key_mem\[2\]\[56\] _06617_ sky130_fd_sc_hd__mux2_2
X_12010_ VGND VPWR _07612_ _07591_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21208_ VGND VPWR _01345_ _06058_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22188_ VGND VPWR VPWR VGND _06578_ _02660_ keymem.key_mem\[2\]\[23\] _06581_ sky130_fd_sc_hd__mux2_2
X_21139_ VGND VPWR _01312_ _06022_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_246_977 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_100_2_Right_172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13961_ VPWR VGND VPWR VGND _09298_ _09245_ _09266_ _09254_ _09433_ sky130_fd_sc_hd__or4_2
XFILLER_0_191_1307 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_57_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12912_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[75\] _08137_ keymem.key_mem\[1\]\[75\]
+ _07901_ _08440_ sky130_fd_sc_hd__a22o_2
X_15700_ VPWR VGND _11156_ keymem.prev_key1_reg\[48\] keymem.prev_key1_reg\[16\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
X_16680_ _02832_ _02834_ _02831_ _02833_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_13892_ VGND VPWR VGND VPWR _09364_ _09291_ _09285_ _09328_ _09306_ sky130_fd_sc_hd__and4_2
XFILLER_0_241_660 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15631_ VPWR VGND VPWR VGND _11080_ _11088_ _11087_ _11077_ _11089_ sky130_fd_sc_hd__or4_2
X_24829_ VGND VPWR VPWR VGND clk _01322_ reset_n keymem.key_mem\[6\]\[54\] sky130_fd_sc_hd__dfrtp_2
X_12843_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[68\] _07667_ keymem.key_mem\[11\]\[68\]
+ _07861_ _08378_ sky130_fd_sc_hd__a22o_2
XFILLER_0_55_1270 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18350_ VPWR VGND _04247_ _04246_ enc_block.round_key\[121\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_68_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15562_ VGND VPWR VGND VPWR _11020_ _10979_ _11021_ _11019_ sky130_fd_sc_hd__nand3_2
XFILLER_0_115_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12774_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[61\] _07595_ keymem.key_mem\[3\]\[61\]
+ _07602_ _08316_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_177_2_Right_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_189_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_90_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14513_ VPWR VGND _09941_ _09982_ _09981_ VPWR VGND sky130_fd_sc_hd__and2_2
X_17301_ VGND VPWR VGND VPWR _11624_ _03395_ _02667_ _02671_ _03397_ sky130_fd_sc_hd__a31o_2
X_11725_ VGND VPWR result[29] _07426_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_138_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15493_ VPWR VGND VGND VPWR _10953_ _10514_ _10562_ sky130_fd_sc_hd__nand2_2
X_18281_ VGND VPWR _04184_ enc_block.block_w1_reg\[18\] _04183_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_51_1167 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_12_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14444_ VPWR VGND VGND VPWR _09440_ _09913_ _09391_ sky130_fd_sc_hd__nor2_2
X_17232_ VGND VPWR _02342_ _03333_ _03335_ _03334_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_37_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_86_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11656_ VPWR VGND VPWR VGND _07391_ aes_core_ctrl_reg\[1\] aes_core_ctrl_reg\[2\]
+ sky130_fd_sc_hd__or2_2
XFILLER_0_126_358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_128_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17163_ VGND VPWR VPWR VGND _03273_ _10735_ _03270_ _03271_ _03272_ sky130_fd_sc_hd__o31a_2
X_14375_ VPWR VGND VPWR VGND _09840_ _09844_ _09841_ _09839_ _09845_ sky130_fd_sc_hd__or4_2
X_16114_ VGND VPWR VGND VPWR _11564_ _11292_ _11565_ _11566_ _11568_ _11567_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_52_665 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13326_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[116\] _07730_ keymem.key_mem\[8\]\[116\]
+ _07541_ _08813_ sky130_fd_sc_hd__a22o_2
XFILLER_0_134_391 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_208_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17094_ VGND VPWR _03211_ _03077_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_12_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_838 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16045_ VPWR VGND VPWR VGND _11405_ _11499_ _11498_ _11293_ _11500_ sky130_fd_sc_hd__or4_2
XFILLER_0_10_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13257_ VGND VPWR enc_block.round_key\[108\] _08751_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_126_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12208_ VGND VPWR _07800_ _07799_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_23_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13188_ VPWR VGND VPWR VGND _08688_ keymem.key_mem\[13\]\[102\] _07588_ keymem.key_mem\[14\]\[102\]
+ _07584_ _08689_ sky130_fd_sc_hd__a221o_2
XFILLER_0_161_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19804_ VGND VPWR _00688_ _05311_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_23_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12139_ VPWR VGND VPWR VGND keymem.key_mem\[4\]\[7\] _07734_ keymem.key_mem\[2\]\[7\]
+ _07733_ _07735_ sky130_fd_sc_hd__a22o_2
X_17996_ VPWR VGND VPWR VGND _03929_ keymem.prev_key1_reg\[122\] sky130_fd_sc_hd__inv_2
XFILLER_0_97_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_252_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19735_ VGND VPWR _00655_ _05275_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16947_ VPWR VGND VPWR VGND _02493_ _02490_ _03078_ key[181] _03077_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_262_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19666_ VGND VPWR VPWR VGND _05227_ _05085_ keymem.key_mem\[12\]\[125\] _05237_ sky130_fd_sc_hd__mux2_2
XFILLER_0_56_1023 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16878_ VGND VPWR VPWR VGND _02986_ keymem.key_mem\[14\]\[46\] _03015_ _03016_ sky130_fd_sc_hd__mux2_2
XFILLER_0_215_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_885 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18617_ VPWR VGND VPWR VGND _04486_ _04459_ _04485_ enc_block.block_w1_reg\[18\]
+ _04424_ _00326_ sky130_fd_sc_hd__a221o_2
XFILLER_0_250_1415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_822 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15829_ VGND VPWR VGND VPWR _11284_ _11278_ _11280_ _11283_ _11285_ sky130_fd_sc_hd__a31o_2
X_19597_ VPWR VGND keymem.key_mem\[12\]\[92\] _05201_ _05094_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_133_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_855 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18548_ VGND VPWR _04424_ _04316_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_133_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18479_ VGND VPWR VGND VPWR _04361_ _03951_ _04362_ _00312_ sky130_fd_sc_hd__a21o_2
XFILLER_0_28_640 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_144_100 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20510_ VGND VPWR _01019_ _05686_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_34_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21490_ VGND VPWR _01478_ _06207_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_55_470 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_846 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20441_ VGND VPWR _05649_ _05533_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23160_ VGND VPWR VGND VPWR _02291_ _07064_ _06888_ keymem.prev_key1_reg\[114\] sky130_fd_sc_hd__o21a_2
XFILLER_0_63_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20372_ VGND VPWR VPWR VGND _05602_ _03252_ keymem.key_mem\[9\]\[71\] _05613_ sky130_fd_sc_hd__mux2_2
XFILLER_0_144_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_139_2_Right_211 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_259_546 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22111_ VGND VPWR VPWR VGND _06538_ _05066_ keymem.key_mem\[3\]\[116\] _06539_ sky130_fd_sc_hd__mux2_2
XFILLER_0_3_773 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_42_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23091_ VGND VPWR VGND VPWR _07021_ _03406_ _06890_ _03408_ _07011_ sky130_fd_sc_hd__a211o_2
XFILLER_0_144_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1096 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_80_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22042_ VPWR VGND keymem.key_mem\[3\]\[83\] _06503_ _06484_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_11_573 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_251_Right_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_140_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_584 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25801_ keymem.prev_key1_reg\[117\] clk _02294_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_242_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23993_ VGND VPWR VPWR VGND clk _00486_ reset_n keymem.key_mem\[13\]\[114\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_242_446 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25732_ keymem.prev_key1_reg\[48\] clk _02225_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22944_ VPWR VGND VPWR VGND _06934_ keymem.prev_key1_reg\[29\] _06926_ sky130_fd_sc_hd__or2_2
XFILLER_0_138_1157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_74_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25663_ VGND VPWR VPWR VGND clk _02156_ reset_n keymem.key_mem\[0\]\[120\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_183_82 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22875_ VGND VPWR _06890_ _10085_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24614_ VGND VPWR VPWR VGND clk _01107_ reset_n keymem.key_mem\[8\]\[95\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_167_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21826_ VGND VPWR VPWR VGND _06377_ _03573_ keymem.key_mem\[4\]\[113\] _06385_ sky130_fd_sc_hd__mux2_2
XFILLER_0_190_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25594_ VGND VPWR VPWR VGND clk _02087_ reset_n keymem.key_mem\[0\]\[51\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_112_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_151_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24545_ VGND VPWR VPWR VGND clk _01038_ reset_n keymem.key_mem\[8\]\[26\] sky130_fd_sc_hd__dfrtp_2
X_21757_ VGND VPWR VPWR VGND _06344_ _03329_ keymem.key_mem\[4\]\[80\] _06349_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_662 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20708_ VGND VPWR VPWR VGND _05783_ _03506_ keymem.key_mem\[8\]\[102\] _05790_ sky130_fd_sc_hd__mux2_2
XFILLER_0_19_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12490_ VPWR VGND VPWR VGND _08058_ keymem.key_mem\[13\]\[34\] _07622_ keymem.key_mem\[8\]\[34\]
+ _07655_ _08059_ sky130_fd_sc_hd__a221o_2
X_24476_ VGND VPWR VPWR VGND clk _00969_ reset_n keymem.key_mem\[9\]\[85\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21688_ VGND VPWR VPWR VGND _06308_ _03024_ keymem.key_mem\[4\]\[47\] _06313_ sky130_fd_sc_hd__mux2_2
XFILLER_0_80_226 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23427_ VGND VPWR VGND VPWR _07295_ _04149_ _07095_ _07296_ enc_block.block_w3_reg\[22\]
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_62_952 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20639_ VGND VPWR VPWR VGND _05747_ _03234_ keymem.key_mem\[8\]\[69\] _05754_ sky130_fd_sc_hd__mux2_2
XFILLER_0_266_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14160_ VGND VPWR VGND VPWR _09629_ keymem.prev_key1_reg\[97\] _09631_ _09589_ sky130_fd_sc_hd__nand3_2
X_23358_ VPWR VGND VPWR VGND _07234_ _07157_ _07232_ sky130_fd_sc_hd__or2_2
XFILLER_0_21_315 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_162_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13111_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[94\] _07742_ keymem.key_mem\[12\]\[94\]
+ _07673_ _08620_ sky130_fd_sc_hd__a22o_2
XFILLER_0_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22309_ VGND VPWR VPWR VGND _06634_ _03339_ keymem.key_mem\[2\]\[81\] _06644_ sky130_fd_sc_hd__mux2_2
X_14091_ VPWR VGND VPWR VGND _09299_ _09317_ _09315_ _09297_ _09562_ sky130_fd_sc_hd__or4_2
X_23289_ VPWR VGND VPWR VGND _07171_ block[8] _04351_ enc_block.block_w1_reg\[8\]
+ _03978_ _07172_ sky130_fd_sc_hd__a221o_2
XFILLER_0_123_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_131_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13042_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[87\] _08449_ _08557_ _08553_ _08558_
+ sky130_fd_sc_hd__o22a_2
X_25028_ VGND VPWR VPWR VGND clk _01521_ reset_n keymem.key_mem\[5\]\[125\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_197_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_123_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17850_ VGND VPWR VPWR VGND _03814_ _03829_ keymem.prev_key0_reg\[75\] _03830_ sky130_fd_sc_hd__mux2_2
XFILLER_0_197_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_219_999 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16801_ VGND VPWR VPWR VGND _02884_ keymem.key_mem\[14\]\[39\] _02945_ _02946_ sky130_fd_sc_hd__mux2_2
XFILLER_0_218_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17781_ VGND VPWR _00194_ _03782_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14993_ VGND VPWR _10457_ _10456_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_101_2_Right_173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19520_ VGND VPWR _00555_ _05160_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16732_ VPWR VGND VPWR VGND _02882_ _02878_ _02876_ key[161] _02875_ _02883_ sky130_fd_sc_hd__a221o_2
X_13944_ VGND VPWR VPWR VGND _09331_ _09246_ _09319_ _09416_ sky130_fd_sc_hd__or3_2
XFILLER_0_202_800 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_191_1148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19451_ VGND VPWR VGND VPWR _05123_ keymem.key_mem_we _02661_ _05121_ _00523_ sky130_fd_sc_hd__a31o_2
X_13875_ VPWR VGND VPWR VGND _09307_ _09291_ _09321_ _09338_ _09347_ sky130_fd_sc_hd__or4_2
XFILLER_0_173_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16663_ VPWR VGND VGND VPWR keymem.prev_key0_reg\[126\] _02816_ _10360_ _02814_ _02815_
+ _02817_ sky130_fd_sc_hd__a311o_2
XFILLER_0_53_1229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18402_ VPWR VGND VPWR VGND _04293_ _04291_ _04290_ enc_block.block_w0_reg\[30\]
+ _03993_ _00304_ sky130_fd_sc_hd__a221o_2
X_15614_ VGND VPWR VPWR VGND _11065_ _11071_ _10493_ _11072_ sky130_fd_sc_hd__or3_2
XFILLER_0_134_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12826_ VPWR VGND VPWR VGND _08362_ keymem.key_mem\[6\]\[66\] _08137_ keymem.key_mem\[8\]\[66\]
+ _07655_ _08363_ sky130_fd_sc_hd__a221o_2
X_19382_ VGND VPWR _00495_ _05082_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16594_ VGND VPWR _02751_ keymem.prev_key0_reg\[59\] keymem.prev_key0_reg\[91\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18333_ VGND VPWR VGND VPWR _02637_ _02612_ _03970_ _04232_ sky130_fd_sc_hd__a21o_2
X_15545_ VPWR VGND VPWR VGND _11003_ _11004_ _10872_ _11002_ sky130_fd_sc_hd__or3b_2
X_12757_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[59\] _08032_ keymem.key_mem\[1\]\[59\]
+ _07799_ _08301_ sky130_fd_sc_hd__a22o_2
XFILLER_0_16_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11708_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[21\] dec_new_block\[21\]
+ _07418_ sky130_fd_sc_hd__mux2_2
XFILLER_0_210_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15476_ VPWR VGND VGND VPWR _10668_ _10936_ _10522_ sky130_fd_sc_hd__nor2_2
X_18264_ VGND VPWR VGND VPWR _11532_ _11502_ _04073_ _04169_ sky130_fd_sc_hd__a21o_2
X_12688_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[52\] _08145_ _08238_ _08234_ _08239_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_71_215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14427_ VPWR VGND VPWR VGND _09891_ _09895_ _09893_ _09889_ _09896_ sky130_fd_sc_hd__or4_2
X_17215_ VGND VPWR VPWR VGND _03020_ keymem.prev_key0_reg\[79\] _03320_ _03319_ _03318_
+ sky130_fd_sc_hd__o211a_2
X_11639_ VPWR VGND VPWR VGND _07378_ keylen sky130_fd_sc_hd__inv_2
X_18195_ VPWR VGND _04106_ _04105_ enc_block.round_key\[107\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_29_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_25_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14358_ VPWR VGND VGND VPWR _09077_ _09828_ _09173_ sky130_fd_sc_hd__nor2_2
XFILLER_0_108_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17146_ key[200] _03258_ keylen _10325_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_180_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13309_ VGND VPWR VGND VPWR _07778_ keymem.key_mem\[3\]\[114\] _08795_ _08797_ _08798_
+ _08736_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_141_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17077_ VGND VPWR VPWR VGND _09710_ _09711_ keymem.prev_key0_reg\[65\] _03196_ sky130_fd_sc_hd__or3_2
X_14289_ VPWR VGND VGND VPWR _09739_ _09746_ _09752_ _09758_ _09759_ sky130_fd_sc_hd__and4b_2
XFILLER_0_64_1369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_668 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_97_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_516 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16028_ VGND VPWR VGND VPWR _11469_ _11482_ _11483_ _11246_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_141_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_196_1037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_23_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_141_1_Left_408 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17979_ VGND VPWR VPWR VGND _03674_ _03917_ keymem.prev_key0_reg\[116\] _03918_ sky130_fd_sc_hd__mux2_2
X_19718_ VGND VPWR _00647_ _05266_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20990_ VGND VPWR _01243_ _05942_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_196_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19649_ VGND VPWR _00616_ _05228_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_149_203 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_149_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22660_ VGND VPWR _02054_ _06801_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_215_1376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_370 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_153_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21611_ VGND VPWR _01534_ _06272_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_36_908 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22591_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[103\] _06775_ _06774_ _05039_ _02011_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_5_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24330_ VGND VPWR VPWR VGND clk _00823_ reset_n keymem.key_mem\[10\]\[67\] sky130_fd_sc_hd__dfrtp_2
X_21542_ VGND VPWR VPWR VGND _06231_ _03538_ keymem.key_mem\[5\]\[107\] _06235_ sky130_fd_sc_hd__mux2_2
XFILLER_0_62_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_69_1225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_941 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24261_ VGND VPWR VPWR VGND clk _00754_ reset_n keymem.key_mem\[11\]\[126\] sky130_fd_sc_hd__dfrtp_2
X_21473_ VPWR VGND VGND VPWR _06199_ keymem.key_mem\[5\]\[74\] _06114_ sky130_fd_sc_hd__nand2_2
XFILLER_0_172_272 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23212_ VPWR VGND VGND VPWR _07102_ _07097_ _07100_ sky130_fd_sc_hd__nand2_2
X_20424_ VGND VPWR _00979_ _05640_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_31_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_86_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24192_ VGND VPWR VPWR VGND clk _00685_ reset_n keymem.key_mem\[11\]\[57\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_261_1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_120_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23143_ VGND VPWR VPWR VGND _07054_ _07053_ keymem.prev_key1_reg\[107\] _07055_ sky130_fd_sc_hd__mux2_2
X_20355_ VGND VPWR _00946_ _05604_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_219_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23074_ VGND VPWR VGND VPWR _07012_ _03336_ _03335_ _03338_ _07011_ sky130_fd_sc_hd__a211o_2
XFILLER_0_140_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20286_ VGND VPWR VPWR VGND _05558_ _02839_ keymem.key_mem\[9\]\[30\] _05568_ sky130_fd_sc_hd__mux2_2
XFILLER_0_80_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1224 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22025_ VGND VPWR VPWR VGND _01727_ _06406_ _03286_ _08922_ _06493_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_216_914 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_216_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_947 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_264_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23976_ VGND VPWR VPWR VGND clk _00469_ reset_n keymem.key_mem\[13\]\[97\] sky130_fd_sc_hd__dfrtp_2
X_11990_ VGND VPWR _07593_ _07592_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_166_2_Left_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22927_ VGND VPWR _02200_ _06922_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25715_ keymem.prev_key1_reg\[31\] clk _02208_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_195_320 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13660_ VGND VPWR _09132_ _08999_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_85_318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25646_ VGND VPWR VPWR VGND clk _02139_ reset_n keymem.key_mem\[0\]\[103\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22858_ VPWR VGND VGND VPWR _03727_ _06877_ _08929_ sky130_fd_sc_hd__nor2_2
XFILLER_0_116_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12611_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[45\] _07778_ keymem.key_mem\[8\]\[45\]
+ _07753_ _08169_ sky130_fd_sc_hd__a22o_2
X_21809_ VGND VPWR VPWR VGND _06366_ _03525_ keymem.key_mem\[4\]\[105\] _06376_ sky130_fd_sc_hd__mux2_2
XFILLER_0_13_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13591_ VGND VPWR VGND VPWR _09063_ _09061_ _09060_ _09047_ _09062_ _09059_ sky130_fd_sc_hd__a32o_2
X_25577_ VGND VPWR VPWR VGND clk _02070_ reset_n keymem.key_mem\[0\]\[34\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_155_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22789_ VGND VPWR _02129_ _06855_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15330_ VPWR VGND VGND VPWR _10792_ _10790_ _10791_ sky130_fd_sc_hd__nand2_2
XFILLER_0_87_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12542_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[39\] _07894_ keymem.key_mem\[8\]\[39\]
+ _07958_ _08106_ sky130_fd_sc_hd__a22o_2
X_24528_ VGND VPWR VPWR VGND clk _01021_ reset_n keymem.key_mem\[8\]\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_727 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_384 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_481 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15261_ VPWR VGND VPWR VGND _10723_ _10724_ _10721_ _10722_ sky130_fd_sc_hd__or3b_2
XFILLER_0_87_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_248 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12473_ VGND VPWR VGND VPWR _08044_ _08008_ keymem.key_mem\[2\]\[32\] _08041_ _08043_
+ sky130_fd_sc_hd__a211o_2
X_24459_ VGND VPWR VPWR VGND clk _00952_ reset_n keymem.key_mem\[9\]\[68\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_34_440 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14212_ VPWR VGND VPWR VGND _09031_ _09065_ _09017_ _09009_ _09683_ sky130_fd_sc_hd__or4_2
X_17000_ VGND VPWR VGND VPWR _02736_ _02735_ _03126_ _03124_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_22_613 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15192_ VPWR VGND VGND VPWR _10655_ _10656_ _10386_ sky130_fd_sc_hd__nor2_2
XFILLER_0_61_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14143_ VGND VPWR VGND VPWR _09294_ _09408_ _09388_ _09443_ _09614_ sky130_fd_sc_hd__o22a_2
XFILLER_0_104_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18951_ VPWR VGND _04787_ _04786_ enc_block.round_key\[52\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_14074_ VPWR VGND _09545_ keymem.prev_key1_reg\[33\] keymem.prev_key1_reg\[1\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_162_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13025_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[86\] _07659_ keymem.key_mem\[10\]\[86\]
+ _08193_ _08542_ sky130_fd_sc_hd__a22o_2
X_17902_ VPWR VGND VGND VPWR _03731_ _03866_ _03424_ sky130_fd_sc_hd__nor2_2
XFILLER_0_238_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18882_ VPWR VGND _04725_ _04724_ enc_block.round_key\[45\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_20_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_219_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_24_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_262 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_158_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17833_ VGND VPWR _03818_ _10371_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_238_96 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_94_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_2_Left_569 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_98_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_83_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17764_ VGND VPWR VPWR VGND _03763_ _03011_ keymem.prev_key0_reg\[46\] _03773_ sky130_fd_sc_hd__mux2_2
X_14976_ VGND VPWR _10440_ _10403_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_102_2_Right_174 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_234_1218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19503_ VGND VPWR _05151_ _05091_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_221_416 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_178_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16715_ VGND VPWR _02866_ key[32] _02867_ _09988_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_13927_ VGND VPWR _09399_ _09398_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_53_1004 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_107_67 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17695_ VGND VPWR _00164_ _03726_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_16_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19434_ VPWR VGND keymem.key_mem\[12\]\[16\] _05114_ _05102_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_76_318 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16646_ VGND VPWR VPWR VGND _02799_ _02800_ keymem.prev_key1_reg\[125\] _02801_ sky130_fd_sc_hd__or3_2
X_13858_ VGND VPWR _09330_ _09329_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_134_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12809_ VPWR VGND VPWR VGND _08347_ keymem.key_mem\[13\]\[64\] _07835_ keymem.key_mem\[2\]\[64\]
+ _07648_ _08348_ sky130_fd_sc_hd__a221o_2
X_19365_ VPWR VGND keymem.key_mem_we _05071_ _03607_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_31_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16577_ VGND VPWR VPWR VGND _02733_ _02734_ keymem.prev_key1_reg\[90\] _02735_ sky130_fd_sc_hd__or3_2
X_13789_ VGND VPWR _09261_ _09260_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_35_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_146_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18316_ VPWR VGND VGND VPWR _04216_ enc_block.block_w2_reg\[13\] enc_block.block_w2_reg\[14\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_225_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15528_ VPWR VGND VPWR VGND _10986_ _10987_ _10523_ _10984_ sky130_fd_sc_hd__or3b_2
XFILLER_0_70_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19296_ VPWR VGND keymem.key_mem_we _05024_ _03466_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_267_1049 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_749 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_169_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_824 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18247_ VGND VPWR _04153_ enc_block.block_w3_reg\[0\] _04152_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15459_ VGND VPWR VGND VPWR _10488_ _10490_ _10919_ _10462_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_5_835 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_154_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18178_ VGND VPWR _04090_ enc_block.block_w1_reg\[18\] _04089_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_128_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_356 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_102_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17129_ VPWR VGND VGND VPWR _03243_ key[198] _10967_ sky130_fd_sc_hd__nand2_2
XFILLER_0_25_1117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_64_1177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_141_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20140_ VGND VPWR _00846_ _05489_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_102_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20071_ VGND VPWR _00813_ _05453_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_176_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_755 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23830_ VGND VPWR VPWR VGND clk _00323_ reset_n enc_block.block_w1_reg\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_256_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_917 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_574 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_164_40 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23761_ keymem.prev_key0_reg\[117\] clk _00258_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20973_ VGND VPWR VGND VPWR _05933_ keymem.key_mem_we _03460_ _05916_ _01235_ sky130_fd_sc_hd__a31o_2
X_22712_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[50\] _06820_ _06819_ _04955_ _02086_
+ sky130_fd_sc_hd__a22o_2
X_25500_ VGND VPWR VPWR VGND clk _01993_ reset_n keymem.key_mem\[1\]\[85\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_73_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_250_1031 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_113_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23692_ keymem.prev_key0_reg\[48\] clk _00189_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_152_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_211_1015 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25431_ VGND VPWR VPWR VGND clk _01924_ reset_n keymem.key_mem\[1\]\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_215_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22643_ VGND VPWR VPWR VGND _06785_ keymem.key_mem\[0\]\[10\] _10836_ _06793_ sky130_fd_sc_hd__mux2_2
XFILLER_0_113_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_211_1059 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_187_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25362_ VGND VPWR VPWR VGND clk _01855_ reset_n keymem.key_mem\[2\]\[75\] sky130_fd_sc_hd__dfrtp_2
X_22574_ VGND VPWR _01999_ _06770_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_187_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24313_ VGND VPWR VPWR VGND clk _00806_ reset_n keymem.key_mem\[10\]\[50\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_8_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21525_ VGND VPWR VPWR VGND _06220_ _03485_ keymem.key_mem\[5\]\[99\] _06226_ sky130_fd_sc_hd__mux2_2
X_25293_ VGND VPWR VPWR VGND clk _01786_ reset_n keymem.key_mem\[2\]\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_111_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_90_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_263_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_16_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_771 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24244_ VGND VPWR VPWR VGND clk _00737_ reset_n keymem.key_mem\[11\]\[109\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_50_218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21456_ VGND VPWR VPWR VGND _06184_ _03209_ keymem.key_mem\[5\]\[66\] _06190_ sky130_fd_sc_hd__mux2_2
XFILLER_0_263_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20407_ VGND VPWR _00971_ _05631_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_160_275 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24175_ VGND VPWR VPWR VGND clk _00668_ reset_n keymem.key_mem\[11\]\[40\] sky130_fd_sc_hd__dfrtp_2
X_21387_ VGND VPWR VPWR VGND _06151_ _02883_ keymem.key_mem\[5\]\[33\] _06154_ sky130_fd_sc_hd__mux2_2
XFILLER_0_32_999 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_248_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1171 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23126_ VGND VPWR VGND VPWR _03502_ _06928_ _03505_ _07043_ sky130_fd_sc_hd__a21o_2
XFILLER_0_113_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20338_ VGND VPWR _00938_ _05595_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_120_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_806 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_60_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23057_ VGND VPWR VGND VPWR _03281_ key[203] _10908_ _07001_ sky130_fd_sc_hd__a21o_2
X_20269_ VGND VPWR _00905_ _05559_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22008_ VPWR VGND keymem.key_mem\[3\]\[67\] _06485_ _06484_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_194_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_44 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_200_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14830_ VGND VPWR VGND VPWR _09411_ _09327_ _09358_ _09450_ _10295_ sky130_fd_sc_hd__a31o_2
XFILLER_0_243_552 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_235_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_208_77 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_215_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_235_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_287 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_8_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14761_ VGND VPWR VGND VPWR _10223_ _09181_ _10224_ _10225_ _10227_ _10226_ sky130_fd_sc_hd__a2111o_2
X_11973_ VPWR VGND VGND VPWR _07531_ _07576_ _07527_ sky130_fd_sc_hd__nor2_2
X_23959_ VGND VPWR VPWR VGND clk _00452_ reset_n keymem.key_mem\[13\]\[80\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_203_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_231_769 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16500_ VGND VPWR _02661_ _02660_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_58_318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13712_ VPWR VGND VGND VPWR _09058_ _09184_ _08958_ sky130_fd_sc_hd__nor2_2
X_14692_ VGND VPWR VGND VPWR _09217_ _09050_ _09102_ _09068_ _10159_ sky130_fd_sc_hd__o22a_2
X_17480_ VGND VPWR VPWR VGND _11092_ _10735_ _03554_ _10328_ _03553_ sky130_fd_sc_hd__o211a_2
XFILLER_0_224_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_131_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16431_ VPWR VGND VPWR VGND _02593_ keymem.prev_key0_reg\[22\] sky130_fd_sc_hd__inv_2
X_13643_ VPWR VGND VPWR VGND _09010_ _09065_ _08971_ _08958_ _09115_ sky130_fd_sc_hd__or4_2
X_25629_ VGND VPWR VPWR VGND clk _02122_ reset_n keymem.key_mem\[0\]\[86\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_131_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19150_ VGND VPWR _00411_ _04934_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16362_ VGND VPWR VGND VPWR _02525_ _11392_ _11230_ _02374_ _02524_ sky130_fd_sc_hd__a211o_2
X_13574_ VGND VPWR VGND VPWR _09046_ _09015_ _09045_ _09044_ _09043_ sky130_fd_sc_hd__and4_2
XFILLER_0_13_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18101_ VPWR VGND VGND VPWR _04019_ _04020_ _03993_ sky130_fd_sc_hd__nor2_2
X_15313_ VGND VPWR VGND VPWR _10775_ _10774_ _10768_ _10759_ _10756_ sky130_fd_sc_hd__and4_2
X_12525_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[37\] _07610_ keymem.key_mem\[11\]\[37\]
+ _08090_ _08091_ sky130_fd_sc_hd__a22o_2
X_16293_ VPWR VGND VPWR VGND _02449_ _02456_ _02454_ _02444_ _02457_ sky130_fd_sc_hd__or4_2
X_19081_ VPWR VGND VGND VPWR _10913_ _04894_ _08921_ sky130_fd_sc_hd__nor2_2
XFILLER_0_240_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18032_ VGND VPWR _03954_ _03953_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_81_376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15244_ VPWR VGND VGND VPWR _10707_ _10705_ _10706_ sky130_fd_sc_hd__nand2_2
X_12456_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[31\] _07683_ keymem.key_mem\[2\]\[31\]
+ _07546_ _08028_ sky130_fd_sc_hd__a22o_2
XFILLER_0_242_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1199 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15175_ VGND VPWR _10639_ _10594_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_23_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12387_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[25\] _07631_ keymem.key_mem\[4\]\[25\]
+ _07913_ _07965_ sky130_fd_sc_hd__a22o_2
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14126_ VPWR VGND VPWR VGND _09595_ _09596_ _09597_ _09593_ _09594_ sky130_fd_sc_hd__or4b_2
XFILLER_0_10_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_266_633 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19983_ VGND VPWR _00771_ _05407_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18934_ VGND VPWR _04771_ enc_block.block_w3_reg\[18\] _04770_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_14057_ VGND VPWR VGND VPWR _09527_ _09526_ _09528_ _09529_ sky130_fd_sc_hd__a21o_2
XFILLER_0_24_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_839 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13008_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[84\] _07725_ keymem.key_mem\[9\]\[84\]
+ _07672_ _08527_ sky130_fd_sc_hd__a22o_2
XFILLER_0_118_11 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18865_ VGND VPWR _04709_ _04600_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_98_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17816_ VGND VPWR _03200_ _09632_ _03806_ _03789_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_175_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_98_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18796_ VGND VPWR _04647_ enc_block.block_w2_reg\[28\] enc_block.block_w0_reg\[13\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_234_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17747_ VGND VPWR _00180_ _03762_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14959_ VPWR VGND VPWR VGND _10423_ enc_block.block_w0_reg\[13\] _08951_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_103_2_Right_175 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17678_ VGND VPWR VGND VPWR _11550_ keymem.prev_key1_reg\[18\] _03715_ _03670_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_134_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19417_ VPWR VGND keymem.key_mem\[12\]\[8\] _05105_ _05102_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_186_161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16629_ VPWR VGND VPWR VGND _02785_ _10325_ _02782_ _02783_ _02784_ _10281_ sky130_fd_sc_hd__o311a_2
XFILLER_0_174_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19348_ VGND VPWR _00484_ _05059_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_84_170 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_169_1245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_2_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19279_ VGND VPWR _00460_ _05014_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_150_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_579 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_72_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1280 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21310_ VGND VPWR _01394_ _06111_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22290_ VGND VPWR _06634_ _06552_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_206_1106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_142_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21241_ VGND VPWR _01361_ _06075_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21172_ VGND VPWR _01328_ _06039_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_106_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_245_806 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20123_ VGND VPWR _00838_ _05480_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_106_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20054_ VGND VPWR _00805_ _05444_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24931_ VGND VPWR VPWR VGND clk _01424_ reset_n keymem.key_mem\[5\]\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24862_ VGND VPWR VPWR VGND clk _01355_ reset_n keymem.key_mem\[6\]\[87\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_198_916 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_213_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_77_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23813_ VGND VPWR VPWR VGND clk _00306_ reset_n enc_block.sword_ctr_reg\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_252_1137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24793_ VGND VPWR VPWR VGND clk _01286_ reset_n keymem.key_mem\[6\]\[18\] sky130_fd_sc_hd__dfrtp_2
X_23744_ keymem.prev_key0_reg\[100\] clk _00241_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20956_ VPWR VGND keymem.key_mem\[7\]\[87\] _05925_ _05899_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_49_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_67_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_113_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23675_ keymem.prev_key0_reg\[31\] clk _00172_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20887_ VGND VPWR VGND VPWR _05888_ keymem.key_mem_we _03091_ _05864_ _01194_ sky130_fd_sc_hd__a31o_2
XFILLER_0_64_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25414_ VGND VPWR VPWR VGND clk _01907_ reset_n keymem.key_mem\[2\]\[127\] sky130_fd_sc_hd__dfrtp_2
X_22626_ VGND VPWR VPWR VGND _06779_ keymem.key_mem\[0\]\[3\] _09992_ _06783_ sky130_fd_sc_hd__mux2_2
XFILLER_0_10_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25345_ VGND VPWR VPWR VGND clk _01838_ reset_n keymem.key_mem\[2\]\[58\] sky130_fd_sc_hd__dfrtp_2
X_22557_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[81\] _06754_ _06753_ _05002_ _01989_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_183_1209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_579 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_51_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_192_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12310_ VGND VPWR _07894_ _07673_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_1_1074 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21508_ VGND VPWR VPWR VGND _06209_ _03426_ keymem.key_mem\[5\]\[91\] _06217_ sky130_fd_sc_hd__mux2_2
X_25276_ VGND VPWR VPWR VGND clk _01769_ reset_n keymem.key_mem\[3\]\[117\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_210_23 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13290_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[112\] _07760_ keymem.key_mem\[1\]\[112\]
+ _07558_ _08781_ sky130_fd_sc_hd__a22o_2
XFILLER_0_84_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22488_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[40\] _06707_ _06706_ _04935_ _01948_
+ sky130_fd_sc_hd__a22o_2
X_24227_ VGND VPWR VPWR VGND clk _00720_ reset_n keymem.key_mem\[11\]\[92\] sky130_fd_sc_hd__dfrtp_2
X_12241_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[13\] _07534_ _07830_ _07826_ _07831_
+ sky130_fd_sc_hd__o22a_2
X_21439_ VGND VPWR VPWR VGND _06173_ _03129_ keymem.key_mem\[5\]\[58\] _06181_ sky130_fd_sc_hd__mux2_2
XFILLER_0_31_240 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24158_ VGND VPWR VPWR VGND clk _00651_ reset_n keymem.key_mem\[11\]\[23\] sky130_fd_sc_hd__dfrtp_2
X_12172_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[9\] _07667_ keymem.key_mem\[8\]\[9\]
+ _07752_ _07766_ sky130_fd_sc_hd__a22o_2
XFILLER_0_124_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_655 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23109_ VGND VPWR VPWR VGND _07032_ _07031_ keymem.prev_key1_reg\[95\] _07033_ sky130_fd_sc_hd__mux2_2
XFILLER_0_21_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24089_ VGND VPWR VPWR VGND clk _00582_ reset_n keymem.key_mem\[12\]\[82\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_198_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16980_ VGND VPWR VGND VPWR _03108_ _11151_ key[184] _03103_ _03107_ sky130_fd_sc_hd__a211o_2
XFILLER_0_124_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15931_ VGND VPWR VGND VPWR _11320_ _11306_ _11253_ _11387_ sky130_fd_sc_hd__a21o_2
XFILLER_0_21_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_159_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18650_ VGND VPWR _04516_ enc_block.block_w3_reg\[13\] enc_block.block_w3_reg\[14\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15862_ VGND VPWR _11318_ _11317_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_64_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17601_ VPWR VGND VGND VPWR _10287_ _03659_ key[254] sky130_fd_sc_hd__nor2_2
XFILLER_0_95_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14813_ VPWR VGND VGND VPWR _10279_ key[134] _10278_ sky130_fd_sc_hd__nand2_2
X_18581_ VPWR VGND VGND VPWR _04454_ _04307_ _04453_ sky130_fd_sc_hd__nand2_2
X_15793_ VPWR VGND VPWR VGND _11172_ _11248_ _11247_ _11166_ _11249_ sky130_fd_sc_hd__or4_2
XFILLER_0_203_235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_231_555 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_157_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_8_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17532_ VGND VPWR VGND VPWR _03599_ _03596_ _03595_ _09637_ _03598_ _09931_ sky130_fd_sc_hd__a32o_2
X_14744_ VGND VPWR VPWR VGND _09173_ _09121_ _09040_ _10210_ sky130_fd_sc_hd__or3_2
XFILLER_0_93_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_98_284 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11956_ VPWR VGND VGND VPWR _07537_ _07559_ _07543_ sky130_fd_sc_hd__nor2_2
XFILLER_0_131_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17463_ VGND VPWR _00119_ _03539_ VPWR VGND sky130_fd_sc_hd__buf_1
X_11887_ VGND VPWR result[110] _07507_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14675_ VPWR VGND _10142_ _10141_ keymem.prev_key1_reg\[101\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_233_1092 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_73_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19202_ VGND VPWR VGND VPWR _04967_ keymem.key_mem_we _03130_ _04924_ _00430_ sky130_fd_sc_hd__a31o_2
X_16414_ VPWR VGND VGND VPWR _11217_ _11238_ _02576_ _11419_ _11302_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_39_362 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13626_ VGND VPWR VPWR VGND _09031_ _08971_ _08957_ _09098_ sky130_fd_sc_hd__or3_2
X_17394_ VGND VPWR VGND VPWR _03152_ key[226] _03479_ _03480_ sky130_fd_sc_hd__a21o_2
XFILLER_0_32_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19133_ VGND VPWR _00405_ _04923_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_166_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16345_ VGND VPWR VGND VPWR _11307_ _11282_ _11369_ _11275_ _11258_ _02508_ sky130_fd_sc_hd__o32a_2
X_13557_ VGND VPWR _09029_ _09028_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_67_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_294 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_150_1_Left_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12508_ VGND VPWR enc_block.round_key\[35\] _08075_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19064_ VGND VPWR VGND VPWR _04884_ keymem.key_mem_we _09992_ _04878_ _00375_ sky130_fd_sc_hd__a31o_2
X_16276_ _11340_ _02440_ _11477_ _11417_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_13488_ enc_block.sword_ctr_reg\[1\] _08960_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[3\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_246_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18015_ VGND VPWR _07375_ enc_block.round\[0\] _03942_ _07374_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_15227_ VPWR VGND VGND VPWR _10618_ _10690_ _10519_ sky130_fd_sc_hd__nor2_2
X_12439_ VPWR VGND VPWR VGND _08012_ keymem.key_mem\[11\]\[29\] _08011_ keymem.key_mem\[4\]\[29\]
+ _07854_ _08013_ sky130_fd_sc_hd__a221o_2
XFILLER_0_246_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15158_ VPWR VGND VGND VPWR _10612_ _10622_ _10519_ sky130_fd_sc_hd__nor2_2
XFILLER_0_267_953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_266_430 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_107_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14109_ VPWR VGND VGND VPWR _09422_ _09580_ _09348_ sky130_fd_sc_hd__nor2_2
X_15089_ VPWR VGND VGND VPWR _10473_ _10553_ _10514_ sky130_fd_sc_hd__nor2_2
X_19966_ VGND VPWR VPWR VGND _05389_ _10662_ keymem.key_mem\[10\]\[8\] _05398_ sky130_fd_sc_hd__mux2_2
XFILLER_0_103_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_997 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_266_485 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_177_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18917_ VGND VPWR _04756_ _04684_ _04755_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19897_ VGND VPWR VPWR VGND _05350_ keymem.key_mem\[11\]\[105\] _03525_ _05360_ sky130_fd_sc_hd__mux2_2
XFILLER_0_38_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18848_ VPWR VGND VPWR VGND _04694_ enc_block.block_w1_reg\[1\] enc_block.block_w1_reg\[2\]
+ sky130_fd_sc_hd__or2_2
XFILLER_0_253_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18779_ VGND VPWR VGND VPWR _04631_ _04505_ _04629_ _04630_ _04632_ sky130_fd_sc_hd__a31o_2
XFILLER_0_145_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_253_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20810_ VPWR VGND keymem.key_mem\[7\]\[19\] _05847_ _05844_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_145_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21790_ VGND VPWR _06366_ _06258_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_104_2_Right_176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_114_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20741_ VGND VPWR _01129_ _05807_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_50_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23460_ VGND VPWR _07325_ enc_block.round_key\[26\] _07324_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20672_ VGND VPWR VPWR VGND _05761_ _03374_ keymem.key_mem\[8\]\[85\] _05771_ sky130_fd_sc_hd__mux2_2
XFILLER_0_174_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22411_ VGND VPWR VPWR VGND _06696_ keymem.key_mem\[1\]\[1\] _09725_ _06698_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_82_1_Left_349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_184_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23391_ VGND VPWR _07263_ _04179_ _02323_ _07096_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_11_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25130_ VGND VPWR VPWR VGND clk _01623_ reset_n keymem.key_mem\[4\]\[99\] sky130_fd_sc_hd__dfrtp_2
X_22342_ VGND VPWR _01876_ _06661_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_264_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25061_ VGND VPWR VPWR VGND clk _01554_ reset_n keymem.key_mem\[4\]\[30\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_225_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22273_ VGND VPWR _01843_ _06625_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_175_2_Left_646 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_130_234 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24012_ VGND VPWR VPWR VGND clk _00505_ reset_n keymem.key_mem\[12\]\[5\] sky130_fd_sc_hd__dfrtp_2
X_21224_ VGND VPWR VPWR VGND _06065_ _03374_ keymem.key_mem\[6\]\[85\] _06067_ sky130_fd_sc_hd__mux2_2
X_21155_ VGND VPWR VPWR VGND _06029_ _03075_ keymem.key_mem\[6\]\[52\] _06031_ sky130_fd_sc_hd__mux2_2
XFILLER_0_121_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20106_ VPWR VGND VGND VPWR _05472_ keymem.key_mem\[10\]\[74\] _05402_ sky130_fd_sc_hd__nand2_2
X_21086_ VGND VPWR _01287_ _05994_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_201_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20037_ VGND VPWR VPWR VGND _05435_ _02964_ keymem.key_mem\[10\]\[41\] _05436_ sky130_fd_sc_hd__mux2_2
X_24914_ VGND VPWR VPWR VGND clk _01407_ reset_n keymem.key_mem\[5\]\[11\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24845_ VGND VPWR VPWR VGND clk _01338_ reset_n keymem.key_mem\[6\]\[70\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_225_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_1149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11810_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[8\] dec_new_block\[72\]
+ _07469_ sky130_fd_sc_hd__mux2_2
X_12790_ VGND VPWR VGND VPWR _07542_ keymem.key_mem\[8\]\[62\] _08326_ _08328_ _08331_
+ _08330_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_241_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21988_ VPWR VGND keymem.key_mem\[3\]\[58\] _06474_ _06469_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_197_267 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24776_ VGND VPWR VPWR VGND clk _01269_ reset_n keymem.key_mem\[6\]\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_157_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_150_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_150_1_Right_751 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11741_ VGND VPWR result[37] _07434_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_138_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23727_ keymem.prev_key0_reg\[83\] clk _00224_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20939_ VGND VPWR _05916_ _05820_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_37_800 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_90_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_165_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14460_ VGND VPWR VPWR VGND _09928_ _09867_ _09870_ _09929_ sky130_fd_sc_hd__mux2_2
X_11672_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[3\] dec_new_block\[3\]
+ _07400_ sky130_fd_sc_hd__mux2_2
XFILLER_0_48_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23658_ keymem.prev_key0_reg\[14\] clk _00155_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_64_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13411_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[124\] _07702_ keymem.key_mem\[2\]\[124\]
+ _07646_ _08890_ sky130_fd_sc_hd__a22o_2
XFILLER_0_3_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14391_ VPWR VGND VPWR VGND _09860_ _09638_ _09794_ key[130] _09544_ _09861_ sky130_fd_sc_hd__a221o_2
X_22609_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[119\] _06777_ _06776_ _05073_ _02027_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_187_1153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_37_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23589_ VGND VPWR VPWR VGND clk _00090_ reset_n keymem.key_mem\[14\]\[78\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_153_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_64_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16130_ VGND VPWR VGND VPWR _11205_ _11380_ _11284_ _11314_ _11584_ sky130_fd_sc_hd__o22a_2
XPHY_EDGE_ROW_265_Right_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13342_ VPWR VGND VPWR VGND _08827_ keymem.key_mem\[5\]\[117\] _08052_ keymem.key_mem\[14\]\[117\]
+ _07963_ _08828_ sky130_fd_sc_hd__a221o_2
XFILLER_0_88_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25328_ VGND VPWR VPWR VGND clk _01821_ reset_n keymem.key_mem\[2\]\[41\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_106_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16061_ VGND VPWR VPWR VGND _11227_ _11289_ _11288_ _11516_ sky130_fd_sc_hd__or3_2
X_13273_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[110\] _07703_ keymem.key_mem\[2\]\[110\]
+ _07647_ _08766_ sky130_fd_sc_hd__a22o_2
XFILLER_0_49_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25259_ VGND VPWR VPWR VGND clk _01752_ reset_n keymem.key_mem\[3\]\[100\] sky130_fd_sc_hd__dfrtp_2
X_15012_ VGND VPWR _10476_ _10469_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12224_ VGND VPWR VGND VPWR _07808_ keymem.key_mem\[12\]\[12\] _07810_ _07814_ _07815_
+ _07663_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_161_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_249_953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_121_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19820_ VPWR VGND VGND VPWR _05320_ keymem.key_mem\[11\]\[68\] _05243_ sky130_fd_sc_hd__nand2_2
X_12155_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[7\] _07645_ _07750_ _07736_ _07751_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_235_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_202_1367 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19751_ VGND VPWR VPWR VGND _05281_ keymem.key_mem\[11\]\[35\] _02904_ _05284_ sky130_fd_sc_hd__mux2_2
XFILLER_0_159_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16963_ VGND VPWR _00066_ _03092_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12086_ VGND VPWR _07685_ _07582_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18702_ VGND VPWR _04562_ _04496_ _04561_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15914_ VGND VPWR _11370_ _11369_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_246_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19682_ VGND VPWR VPWR VGND _05247_ keymem.key_mem\[11\]\[2\] _09862_ _05248_ sky130_fd_sc_hd__mux2_2
X_16894_ VGND VPWR _09513_ key[48] _03030_ _03029_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_194_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18633_ VPWR VGND VPWR VGND _04500_ block[84] _04487_ enc_block.block_w2_reg\[20\]
+ _04425_ _04501_ sky130_fd_sc_hd__a221o_2
XFILLER_0_246_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15845_ VPWR VGND VGND VPWR _11300_ _11301_ _11255_ sky130_fd_sc_hd__nor2_2
XFILLER_0_204_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_182_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18564_ _04437_ _04439_ _04065_ _04438_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_91_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15776_ VGND VPWR VGND VPWR _11232_ _11165_ _11164_ keymem.prev_key1_reg\[18\] _08955_
+ _08942_ sky130_fd_sc_hd__a32o_2
XFILLER_0_59_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12988_ VPWR VGND VPWR VGND _08508_ keymem.key_mem\[14\]\[82\] _07782_ keymem.key_mem\[2\]\[82\]
+ _08116_ _08509_ sky130_fd_sc_hd__a221o_2
XFILLER_0_86_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_235_1198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17515_ VPWR VGND _09533_ _03584_ _03583_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_172_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14727_ VGND VPWR _10194_ _10193_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18495_ _04375_ _04377_ _04294_ _04376_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_11939_ VGND VPWR _07542_ _07541_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_24_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17446_ VPWR VGND VPWR VGND _03524_ _03521_ _03520_ key[233] _03366_ _03525_ sky130_fd_sc_hd__a221o_2
XFILLER_0_138_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14658_ VGND VPWR VGND VPWR _09333_ _09466_ _09330_ _09475_ _10125_ sky130_fd_sc_hd__o22a_2
X_13609_ VPWR VGND VPWR VGND _09014_ _09015_ _08991_ _09001_ _09081_ sky130_fd_sc_hd__or4_2
X_17377_ VGND VPWR VGND VPWR _03465_ _09637_ _03464_ _03463_ sky130_fd_sc_hd__o21a_2
X_14589_ VPWR VGND VGND VPWR _09420_ _10057_ _09353_ sky130_fd_sc_hd__nor2_2
XFILLER_0_156_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_376 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19116_ VGND VPWR VGND VPWR _04913_ keymem.key_mem_we _02743_ _04908_ _00398_ sky130_fd_sc_hd__a31o_2
XFILLER_0_40_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16328_ _02486_ _02491_ keymem.prev_key1_reg\[85\] _02487_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_232_Right_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19047_ VGND VPWR VGND VPWR _03959_ block[63] _04872_ _04871_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_67_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16259_ VGND VPWR VGND VPWR _02423_ _11400_ _11386_ _11336_ _11246_ _02422_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_28_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_207_1289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_11_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19949_ VGND VPWR _05389_ _05388_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22960_ VGND VPWR _02212_ _06943_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_254_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_156_52 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_173_1208 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_78_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21911_ VPWR VGND keymem.key_mem\[3\]\[22\] _06433_ _06427_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_156_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_257_1390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22891_ VGND VPWR _02186_ _06900_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_39_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21842_ VGND VPWR _01644_ _06393_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24630_ VGND VPWR VPWR VGND clk _01123_ reset_n keymem.key_mem\[8\]\[111\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_190_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24561_ VGND VPWR VPWR VGND clk _01054_ reset_n keymem.key_mem\[8\]\[42\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_210_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21773_ VGND VPWR _01611_ _06357_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_105_2_Right_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_172_95 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20724_ VGND VPWR _01121_ _05798_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23512_ VGND VPWR VPWR VGND clk _00013_ reset_n keymem.key_mem\[14\]\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_147_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_19_833 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24492_ VGND VPWR VPWR VGND clk _00985_ reset_n keymem.key_mem\[9\]\[101\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_188_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23443_ VGND VPWR _07310_ enc_block.round_key\[24\] _07309_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_92_268 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20655_ VGND VPWR _01088_ _05762_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_135_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_18_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23374_ VGND VPWR _07248_ enc_block.block_w3_reg\[25\] enc_block.block_w1_reg\[9\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20586_ VGND VPWR _01055_ _05726_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_184_1359 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1312 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_162_178 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_33_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25113_ VGND VPWR VPWR VGND clk _01606_ reset_n keymem.key_mem\[4\]\[82\] sky130_fd_sc_hd__dfrtp_2
X_22325_ VGND VPWR _01868_ _06652_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_46_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25044_ VGND VPWR VPWR VGND clk _01537_ reset_n keymem.key_mem\[4\]\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_582 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22256_ VGND VPWR _01835_ _06616_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_225_1389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_83_1191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_267_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21207_ VGND VPWR VPWR VGND _06052_ _03306_ keymem.key_mem\[6\]\[77\] _06058_ sky130_fd_sc_hd__mux2_2
XFILLER_0_264_219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22187_ VGND VPWR _01802_ _06580_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_257_260 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21138_ VGND VPWR VPWR VGND _06018_ _02998_ keymem.key_mem\[6\]\[44\] _06022_ sky130_fd_sc_hd__mux2_2
XFILLER_0_233_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13960_ VPWR VGND VGND VPWR _09431_ _09383_ _09432_ _09378_ _09410_ sky130_fd_sc_hd__o22ai_2
X_21069_ VPWR VGND VGND VPWR _05986_ keymem.key_mem\[6\]\[11\] _05985_ sky130_fd_sc_hd__nand2_2
XFILLER_0_96_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12911_ VGND VPWR enc_block.round_key\[74\] _08439_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_236_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13891_ VPWR VGND VGND VPWR _09362_ _09363_ _09361_ sky130_fd_sc_hd__nor2_2
XFILLER_0_9_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15630_ VPWR VGND VPWR VGND _10760_ _10950_ _10843_ _10763_ _11088_ sky130_fd_sc_hd__or4_2
XFILLER_0_57_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24828_ VGND VPWR VPWR VGND clk _01321_ reset_n keymem.key_mem\[6\]\[53\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_236_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12842_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[68\] _07984_ keymem.key_mem\[2\]\[68\]
+ _07816_ _08377_ sky130_fd_sc_hd__a22o_2
XFILLER_0_9_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_694 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15561_ VGND VPWR VGND VPWR _10184_ _10360_ _11020_ _10168_ sky130_fd_sc_hd__nand3_2
XFILLER_0_55_1282 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12773_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[61\] _07578_ keymem.key_mem\[1\]\[61\]
+ _07557_ _08315_ sky130_fd_sc_hd__a22o_2
X_24759_ VGND VPWR VPWR VGND clk _01252_ reset_n keymem.key_mem\[7\]\[112\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_68_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_1_Right_752 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17300_ VGND VPWR VGND VPWR _02671_ _02667_ _03396_ _03395_ sky130_fd_sc_hd__a21oi_2
X_14512_ VGND VPWR VGND VPWR _09954_ _09981_ _09972_ _09980_ _09966_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_90_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18280_ VPWR VGND _04183_ enc_block.block_w0_reg\[27\] enc_block.block_w1_reg\[23\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_83_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11724_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[29\] dec_new_block\[29\]
+ _07426_ sky130_fd_sc_hd__mux2_2
X_15492_ VPWR VGND VPWR VGND _10951_ _10952_ _10841_ _10950_ sky130_fd_sc_hd__or3b_2
XFILLER_0_83_246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_138_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17231_ VGND VPWR VGND VPWR _11536_ _11535_ _03334_ _03332_ sky130_fd_sc_hd__a21oi_2
X_14443_ VPWR VGND VGND VPWR _09911_ _09910_ _09361_ _09360_ _09553_ _09912_ sky130_fd_sc_hd__a311o_2
X_11655_ VPWR VGND VPWR VGND keymem.ready_new keymem.key_mem_we _07390_ _07366_ keymem.key_mem_ctrl_reg\[0\]
+ _00009_ sky130_fd_sc_hd__a221o_2
XFILLER_0_138_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_167_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17162_ VPWR VGND VPWR VGND _03272_ key[74] _11543_ sky130_fd_sc_hd__or2_2
X_14374_ VPWR VGND VPWR VGND _09842_ _09843_ _09844_ _09219_ _09020_ sky130_fd_sc_hd__or4b_2
XFILLER_0_128_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_243_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16113_ VPWR VGND VGND VPWR _11280_ _11567_ _11336_ sky130_fd_sc_hd__nor2_2
XFILLER_0_247_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13325_ VGND VPWR enc_block.round_key\[115\] _08812_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_52_677 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17093_ VGND VPWR _00078_ _03210_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_51_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_208_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16044_ VGND VPWR VGND VPWR _11385_ _11320_ _11499_ _11329_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_204_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13256_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[108\] _08714_ _08750_ _08746_ _08751_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_0_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12207_ VGND VPWR _07799_ _07624_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13187_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[102\] _07809_ keymem.key_mem\[12\]\[102\]
+ _07807_ _08688_ sky130_fd_sc_hd__a22o_2
XFILLER_0_62_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19803_ VGND VPWR VPWR VGND _05303_ keymem.key_mem\[11\]\[60\] _03150_ _05311_ sky130_fd_sc_hd__mux2_2
XFILLER_0_257_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12138_ VGND VPWR _07734_ _07551_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_264_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17995_ VGND VPWR VGND VPWR _03736_ keymem.prev_key0_reg\[121\] _03928_ _00262_ sky130_fd_sc_hd__a21o_2
X_19734_ VGND VPWR VPWR VGND _05270_ keymem.key_mem\[11\]\[27\] _02765_ _05275_ sky130_fd_sc_hd__mux2_2
X_12069_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[3\] _07668_ keymem.key_mem\[14\]\[3\]
+ _07666_ _07669_ sky130_fd_sc_hd__a22o_2
X_16946_ VGND VPWR _03077_ _09522_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_236_499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19665_ VGND VPWR _00624_ _05236_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16877_ VGND VPWR VGND VPWR _03015_ _03013_ _03010_ _03008_ _03014_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_254_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18616_ VPWR VGND VGND VPWR _04380_ _04486_ _04179_ sky130_fd_sc_hd__nor2_2
X_15828_ VGND VPWR _11284_ _11257_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_255_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19596_ VGND VPWR VGND VPWR _05200_ keymem.key_mem_we _03427_ _05187_ _00591_ sky130_fd_sc_hd__a31o_2
XFILLER_0_205_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_215_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18547_ VPWR VGND VPWR VGND _04423_ _04291_ _04422_ enc_block.block_w1_reg\[11\]
+ _04317_ _00319_ sky130_fd_sc_hd__a221o_2
X_15759_ VPWR VGND VPWR VGND _11215_ enc_block.block_w0_reg\[16\] _08995_ sky130_fd_sc_hd__or2_2
XFILLER_0_133_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_176_259 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_142_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18478_ VGND VPWR VPWR VGND _04316_ enc_block.block_w1_reg\[4\] _04030_ _04362_ sky130_fd_sc_hd__mux2_2
XFILLER_0_47_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_63_909 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_200_580 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_150_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17429_ VGND VPWR VPWR VGND _10327_ key[103] _03510_ _02936_ _10328_ sky130_fd_sc_hd__o211a_2
XFILLER_0_117_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20440_ VGND VPWR _00987_ _05648_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_144_156 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20371_ VGND VPWR _00954_ _05612_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_207_1020 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_207_1031 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22110_ VGND VPWR _06538_ _06402_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23090_ VGND VPWR VGND VPWR _02265_ _07020_ _07010_ keymem.prev_key1_reg\[88\] sky130_fd_sc_hd__o21a_2
XFILLER_0_80_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_247_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22041_ VGND VPWR VGND VPWR _06502_ keymem.key_mem_we _03347_ _06498_ _01734_ sky130_fd_sc_hd__a31o_2
XFILLER_0_144_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25800_ keymem.prev_key1_reg\[116\] clk _02293_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_214_105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23992_ VGND VPWR VPWR VGND clk _00485_ reset_n keymem.key_mem\[13\]\[113\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_1200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_436 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25731_ keymem.prev_key1_reg\[47\] clk _02224_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22943_ VGND VPWR VGND VPWR _02205_ _06933_ _06916_ keymem.prev_key1_reg\[28\] sky130_fd_sc_hd__o21a_2
XFILLER_0_39_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25662_ VGND VPWR VPWR VGND clk _02155_ reset_n keymem.key_mem\[0\]\[119\] sky130_fd_sc_hd__dfrtp_2
X_22874_ VGND VPWR VGND VPWR _06888_ _06887_ _02180_ _06889_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_151_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_223_694 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_183_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24613_ VGND VPWR VPWR VGND clk _01106_ reset_n keymem.key_mem\[8\]\[94\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_91_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21825_ VGND VPWR _01636_ _06384_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25593_ VGND VPWR VPWR VGND clk _02086_ reset_n keymem.key_mem\[0\]\[50\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_167_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21756_ VGND VPWR _01603_ _06348_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24544_ VGND VPWR VPWR VGND clk _01037_ reset_n keymem.key_mem\[8\]\[25\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_52_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_106_2_Right_178 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20707_ VGND VPWR _01113_ _05789_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_65_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21687_ VGND VPWR _01570_ _06312_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24475_ VGND VPWR VPWR VGND clk _00968_ reset_n keymem.key_mem\[9\]\[84\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_1117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_119_2_Left_590 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23426_ VGND VPWR _07295_ enc_block.round_key\[22\] _07294_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20638_ VGND VPWR VGND VPWR _05676_ _03227_ _01080_ _05753_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_184_1167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23357_ VPWR VGND VGND VPWR _07233_ _07157_ _07232_ sky130_fd_sc_hd__nand2_2
X_20569_ VGND VPWR _01047_ _05717_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_150_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_202_Right_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13110_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[94\] _07760_ keymem.key_mem\[4\]\[94\]
+ _08077_ _08619_ sky130_fd_sc_hd__a22o_2
XFILLER_0_260_1033 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22308_ VGND VPWR _01860_ _06643_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14090_ VPWR VGND VGND VPWR _09561_ _09558_ _09560_ sky130_fd_sc_hd__nand2_2
XFILLER_0_162_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23288_ _07169_ _07171_ _03982_ _07170_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_131_384 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13041_ VGND VPWR VGND VPWR _08557_ _07731_ keymem.key_mem\[13\]\[87\] _08554_ _08556_
+ sky130_fd_sc_hd__a211o_2
X_22239_ VGND VPWR _01827_ _06607_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25027_ VGND VPWR VPWR VGND clk _01520_ reset_n keymem.key_mem\[5\]\[124\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_162_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_400 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_138_2_Left_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_245_252 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16800_ VGND VPWR VGND VPWR _02945_ _10838_ key[167] _02939_ _02944_ sky130_fd_sc_hd__a211o_2
XFILLER_0_121_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17780_ VGND VPWR VPWR VGND _03777_ _03781_ keymem.prev_key0_reg\[53\] _03782_ sky130_fd_sc_hd__mux2_2
X_14992_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[13\] _08954_ _10456_ _08941_ _10422_
+ _10423_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_233_425 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16731_ VGND VPWR VPWR VGND _09635_ _02879_ _02882_ _02496_ _02881_ sky130_fd_sc_hd__o211a_2
X_13943_ VGND VPWR _09415_ _09375_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_211_Right_80 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19450_ VPWR VGND keymem.key_mem\[12\]\[23\] _05123_ _05116_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_18_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_2_Right_140 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_72_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16662_ VGND VPWR VGND VPWR _10261_ _10243_ _02816_ _09240_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_242_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13874_ VGND VPWR VGND VPWR _09346_ _09295_ _09248_ _09325_ _09345_ sky130_fd_sc_hd__a211o_2
X_18401_ VPWR VGND VGND VPWR _04292_ _04293_ _03974_ sky130_fd_sc_hd__nor2_2
XFILLER_0_173_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15613_ VPWR VGND VPWR VGND _11068_ _10700_ _11069_ _11070_ _11071_ sky130_fd_sc_hd__or4bb_2
X_12825_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[66\] _07812_ keymem.key_mem\[11\]\[66\]
+ _07658_ _08362_ sky130_fd_sc_hd__a22o_2
X_19381_ VGND VPWR VPWR VGND _05067_ _05081_ keymem.key_mem\[13\]\[123\] _05082_ sky130_fd_sc_hd__mux2_2
XFILLER_0_201_344 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16593_ VGND VPWR _02750_ keymem.prev_key0_reg\[123\] _02749_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18332_ VPWR VGND _04231_ _04230_ enc_block.round_key\[119\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15544_ VGND VPWR VPWR VGND _10469_ _10568_ _10500_ _11003_ sky130_fd_sc_hd__or3_2
XFILLER_0_70_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12756_ VGND VPWR VGND VPWR _07877_ keymem.key_mem\[10\]\[59\] _08299_ _08300_ sky130_fd_sc_hd__a21o_2
XFILLER_0_29_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_152_1_Right_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_56_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_1085 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11707_ VGND VPWR result[20] _07417_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18263_ VPWR VGND _04168_ _04167_ enc_block.round_key\[113\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15475_ VGND VPWR VGND VPWR _10931_ _10934_ _10935_ _10564_ _10932_ sky130_fd_sc_hd__nor4_2
XFILLER_0_38_972 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_25_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12687_ VGND VPWR VGND VPWR _08238_ _08096_ keymem.key_mem\[5\]\[52\] _08235_ _08237_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_210_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17214_ VGND VPWR VGND VPWR _03319_ _09513_ _10732_ key[79] sky130_fd_sc_hd__o21a_2
X_14426_ VPWR VGND VPWR VGND _09579_ _09618_ _09617_ _09894_ _09895_ sky130_fd_sc_hd__or4_2
X_18194_ VPWR VGND VPWR VGND _04104_ block[107] _04076_ enc_block.block_w2_reg\[11\]
+ _04007_ _04105_ sky130_fd_sc_hd__a221o_2
X_11638_ VGND VPWR VPWR VGND _00000_ _07374_ _07377_ _07376_ enc_block.sword_ctr_inc
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_126_167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17145_ VGND VPWR VPWR VGND _03256_ _03257_ keymem.prev_key0_reg\[72\] _10327_ _10655_
+ sky130_fd_sc_hd__a31oi_2
XFILLER_0_141_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14357_ VGND VPWR VGND VPWR _09816_ _09826_ _09827_ _09808_ _09822_ sky130_fd_sc_hd__nor4_2
XFILLER_0_97_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_496 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13308_ VPWR VGND VPWR VGND _08796_ keymem.key_mem\[5\]\[114\] _07683_ keymem.key_mem\[8\]\[114\]
+ _07929_ _08797_ sky130_fd_sc_hd__a221o_2
X_17076_ VGND VPWR _00076_ _03195_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_180_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14288_ VPWR VGND VGND VPWR _09755_ _09361_ _09753_ _09248_ _09758_ _09757_ sky130_fd_sc_hd__o221a_2
XFILLER_0_141_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16027_ VGND VPWR _11482_ _11329_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_23_1001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_256_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13239_ VPWR VGND VPWR VGND _08734_ keymem.key_mem\[9\]\[107\] _07717_ keymem.key_mem\[12\]\[107\]
+ _07621_ _08735_ sky130_fd_sc_hd__a221o_2
XFILLER_0_23_1045 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_196_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17978_ VGND VPWR VPWR VGND _03281_ key[244] keymem.prev_key1_reg\[116\] _03917_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_97_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_1_Left_358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_137_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16929_ VGND VPWR VPWR VGND _09521_ key[179] keymem.prev_key1_reg\[51\] _03062_ sky130_fd_sc_hd__mux2_2
X_19717_ VGND VPWR VPWR VGND _05259_ keymem.key_mem\[11\]\[19\] _02410_ _05266_ sky130_fd_sc_hd__mux2_2
XFILLER_0_224_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1300 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19648_ VGND VPWR VPWR VGND _05227_ _05066_ keymem.key_mem\[12\]\[116\] _05228_ sky130_fd_sc_hd__mux2_2
XFILLER_0_79_349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19579_ VPWR VGND keymem.key_mem\[12\]\[83\] _05192_ _05173_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_220_653 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_184_2_Left_655 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_215_1388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21610_ VGND VPWR VPWR VGND _06263_ _10835_ keymem.key_mem\[4\]\[10\] _06272_ sky130_fd_sc_hd__mux2_2
XFILLER_0_87_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22590_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[102\] _06775_ _06774_ _05037_ _02010_
+ sky130_fd_sc_hd__a22o_2
X_21541_ VGND VPWR _01502_ _06234_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_157_270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_62_216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1448 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_56_791 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_69_1237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24260_ VGND VPWR VPWR VGND clk _00753_ reset_n keymem.key_mem\[11\]\[125\] sky130_fd_sc_hd__dfrtp_2
X_21472_ VGND VPWR _01469_ _06198_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_248_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_430 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_105_318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23211_ VPWR VGND VPWR VGND _07101_ _07097_ _07100_ sky130_fd_sc_hd__or2_2
XFILLER_0_244_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20423_ VGND VPWR VPWR VGND _05638_ _03460_ keymem.key_mem\[9\]\[95\] _05640_ sky130_fd_sc_hd__mux2_2
X_24191_ VGND VPWR VPWR VGND clk _00684_ reset_n keymem.key_mem\[11\]\[56\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_43_496 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_113_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23142_ VGND VPWR _07054_ _06880_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20354_ VGND VPWR VPWR VGND _05602_ _03173_ keymem.key_mem\[9\]\[62\] _05604_ sky130_fd_sc_hd__mux2_2
XFILLER_0_247_517 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23073_ VGND VPWR _07011_ _06883_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_45_1270 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20285_ VGND VPWR _00913_ _05567_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_228_731 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22024_ VPWR VGND VGND VPWR _06493_ keymem.key_mem\[3\]\[75\] _06406_ sky130_fd_sc_hd__nand2_2
XFILLER_0_80_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_937 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_76_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_118_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23975_ VGND VPWR VPWR VGND clk _00468_ reset_n keymem.key_mem\[13\]\[96\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_1030 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25714_ keymem.prev_key1_reg\[30\] clk _02207_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_3_Left_271 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22926_ VGND VPWR VPWR VGND _06914_ _06921_ keymem.prev_key1_reg\[23\] _06922_ sky130_fd_sc_hd__mux2_2
X_25645_ VGND VPWR VPWR VGND clk _02138_ reset_n keymem.key_mem\[0\]\[102\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_190_1171 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_195_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22857_ VGND VPWR VGND VPWR _07383_ keymem.ready keymem.ready_new _02176_ sky130_fd_sc_hd__a21o_2
XFILLER_0_78_382 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12610_ VGND VPWR VGND VPWR _07737_ keymem.key_mem\[1\]\[45\] _08166_ _08167_ _08168_
+ _07574_ sky130_fd_sc_hd__a2111o_2
X_21808_ VGND VPWR _01628_ _06375_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13590_ VGND VPWR VGND VPWR _09062_ _09015_ _08991_ _09044_ _09043_ sky130_fd_sc_hd__and4_2
X_25576_ VGND VPWR VPWR VGND clk _02069_ reset_n keymem.key_mem\[0\]\[33\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22788_ VGND VPWR VPWR VGND _06784_ keymem.key_mem\[0\]\[93\] _03444_ _06855_ sky130_fd_sc_hd__mux2_2
XFILLER_0_210_185 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_151_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_107_2_Right_179 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12541_ VGND VPWR enc_block.round_key\[38\] _08105_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24527_ VGND VPWR VPWR VGND clk _01020_ reset_n keymem.key_mem\[8\]\[8\] sky130_fd_sc_hd__dfrtp_2
X_21739_ VGND VPWR _01595_ _06339_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_4_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15260_ VGND VPWR VGND VPWR _10682_ _10496_ _10520_ _10672_ _10646_ _10723_ sky130_fd_sc_hd__o32a_2
XFILLER_0_227_1204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24458_ VGND VPWR VPWR VGND clk _00951_ reset_n keymem.key_mem\[9\]\[67\] sky130_fd_sc_hd__dfrtp_2
X_12472_ VPWR VGND VPWR VGND _08042_ keymem.key_mem\[5\]\[32\] _07597_ keymem.key_mem\[4\]\[32\]
+ _07552_ _08043_ sky130_fd_sc_hd__a221o_2
XFILLER_0_46_290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_87_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14211_ VGND VPWR VGND VPWR _09091_ _09080_ _09153_ _09102_ _09682_ sky130_fd_sc_hd__o22a_2
XFILLER_0_34_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23409_ VPWR VGND VPWR VGND _07279_ block[20] _04837_ enc_block.block_w0_reg\[20\]
+ _04504_ _07280_ sky130_fd_sc_hd__a221o_2
XFILLER_0_163_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15191_ VGND VPWR _10655_ keymem.prev_key0_reg\[104\] _10654_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_24389_ VGND VPWR VPWR VGND clk _00882_ reset_n keymem.key_mem\[10\]\[126\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_22_636 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14142_ VGND VPWR VGND VPWR _09495_ _09403_ _09444_ _09416_ _09613_ sky130_fd_sc_hd__o22a_2
XFILLER_0_50_956 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_205_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18950_ VPWR VGND VPWR VGND _04785_ block[52] _04744_ enc_block.block_w3_reg\[20\]
+ _04666_ _04786_ sky130_fd_sc_hd__a221o_2
XFILLER_0_123_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14073_ VGND VPWR _09544_ _09543_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_266_837 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_63_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13024_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[86\] _07902_ keymem.key_mem\[4\]\[86\]
+ _07693_ _08541_ sky130_fd_sc_hd__a22o_2
X_17901_ VGND VPWR VGND VPWR _03732_ keymem.prev_key1_reg\[91\] _03864_ _03865_ sky130_fd_sc_hd__a21o_2
X_18881_ VPWR VGND VPWR VGND _04723_ block[45] _04351_ enc_block.block_w0_reg\[13\]
+ _03978_ _04724_ sky130_fd_sc_hd__a221o_2
XFILLER_0_123_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_238_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17832_ VGND VPWR _00210_ _03817_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_246_572 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_94_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_447 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17763_ VGND VPWR _00186_ _03772_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_98_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14975_ VGND VPWR _10439_ _10392_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_238_1366 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19502_ VGND VPWR VGND VPWR _05150_ keymem.key_mem_we _03025_ _05135_ _00547_ sky130_fd_sc_hd__a31o_2
XFILLER_0_254_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16714_ VGND VPWR _02866_ _09512_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13926_ VGND VPWR VPWR VGND _09299_ _09315_ _09319_ _09398_ sky130_fd_sc_hd__or3_2
X_17694_ VGND VPWR VPWR VGND _03723_ _03725_ keymem.prev_key0_reg\[23\] _03726_ sky130_fd_sc_hd__mux2_2
XFILLER_0_107_79 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19433_ VGND VPWR VGND VPWR _05113_ keymem.key_mem_we _11149_ _05109_ _00515_ sky130_fd_sc_hd__a31o_2
XFILLER_0_16_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_69_2_Right_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_134_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_186_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16645_ _11301_ _02800_ keymem.rcon_logic.tmp_rcon\[6\] _02536_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__and3_2
X_13857_ VPWR VGND VPWR VGND _09328_ _09309_ _09285_ _09306_ _09329_ sky130_fd_sc_hd__or4_2
XFILLER_0_173_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12808_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[64\] _07690_ keymem.key_mem\[11\]\[64\]
+ _07809_ _08347_ sky130_fd_sc_hd__a22o_2
X_19364_ VGND VPWR _00489_ _05070_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_186_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16576_ _02724_ _02734_ keymem.prev_key1_reg\[122\] _02725_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_13788_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[26\] _09003_ _09260_ _09255_ _09258_
+ _09259_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_201_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_70_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18315_ VPWR VGND _04215_ _04214_ enc_block.block_w0_reg\[30\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_123_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15527_ VPWR VGND VGND VPWR _10612_ _10608_ _10520_ _10565_ _10986_ _10985_ sky130_fd_sc_hd__o221a_2
X_19295_ VGND VPWR VGND VPWR _05023_ keymem.key_mem_we _03460_ _04999_ _00467_ sky130_fd_sc_hd__a31o_2
X_12739_ VGND VPWR VGND VPWR _08285_ _07901_ keymem.key_mem\[1\]\[57\] _08282_ _08284_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_139_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_32_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_153_1_Right_754 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_57_599 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_84_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_120_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_123_89 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_31_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18246_ VGND VPWR _04152_ enc_block.block_w1_reg\[23\] enc_block.block_w0_reg\[24\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_218_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15458_ VGND VPWR VGND VPWR _10522_ _10543_ _10918_ _10541_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_199_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14409_ VPWR VGND VPWR VGND _09762_ _09877_ _09781_ _09554_ _09878_ sky130_fd_sc_hd__or4_2
XFILLER_0_245_1337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18177_ VGND VPWR _04089_ enc_block.block_w3_reg\[2\] enc_block.block_w0_reg\[26\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_772 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15389_ VPWR VGND VPWR VGND _10763_ _10849_ _10846_ _10626_ _10850_ sky130_fd_sc_hd__or4_2
XFILLER_0_0_1481 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17128_ VGND VPWR VGND VPWR _03242_ _02928_ _02927_ key[70] sky130_fd_sc_hd__o21a_2
XFILLER_0_13_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_145_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_466 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17059_ VGND VPWR VGND VPWR _02855_ _02854_ _03180_ _03178_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_257_848 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_141_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_180_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20070_ VGND VPWR VPWR VGND _05446_ _03119_ keymem.key_mem\[10\]\[57\] _05453_ sky130_fd_sc_hd__mux2_2
XFILLER_0_106_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_141_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_57_84 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_252_553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_213_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23760_ keymem.prev_key0_reg\[116\] clk _00257_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20972_ VPWR VGND keymem.key_mem\[7\]\[95\] _05933_ _05823_ VPWR VGND sky130_fd_sc_hd__and2_2
X_22711_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[49\] _06820_ _06819_ _04953_ _02085_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_152_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23691_ keymem.prev_key0_reg\[47\] clk _00188_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_191_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25430_ VGND VPWR VPWR VGND clk _01923_ reset_n keymem.key_mem\[1\]\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_152_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_211_1027 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22642_ VGND VPWR _02045_ _06792_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_87_190 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_113_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22573_ VGND VPWR VPWR VGND _06701_ keymem.key_mem\[1\]\[91\] _03427_ _06770_ sky130_fd_sc_hd__mux2_2
X_25361_ VGND VPWR VPWR VGND clk _01854_ reset_n keymem.key_mem\[2\]\[74\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_536 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24312_ VGND VPWR VPWR VGND clk _00805_ reset_n keymem.key_mem\[10\]\[49\] sky130_fd_sc_hd__dfrtp_2
X_21524_ VGND VPWR _01494_ _06225_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25292_ VGND VPWR VPWR VGND clk _01785_ reset_n keymem.key_mem\[2\]\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_185_1251 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_146_1202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21455_ VGND VPWR _01461_ _06189_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_263_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24243_ VGND VPWR VPWR VGND clk _00736_ reset_n keymem.key_mem\[11\]\[108\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_307 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20406_ VGND VPWR VPWR VGND _05627_ _03393_ keymem.key_mem\[9\]\[87\] _05631_ sky130_fd_sc_hd__mux2_2
X_24174_ VGND VPWR VPWR VGND clk _00667_ reset_n keymem.key_mem\[11\]\[39\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_181_1148 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21386_ VGND VPWR _01428_ _06153_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_226_1281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_163_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23125_ VGND VPWR _02278_ _07042_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20337_ VGND VPWR VPWR VGND _05591_ _03091_ keymem.key_mem\[9\]\[54\] _05595_ sky130_fd_sc_hd__mux2_2
XFILLER_0_248_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23056_ VGND VPWR VGND VPWR _06881_ _03276_ _02251_ _07000_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_21_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_120_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20268_ VGND VPWR VPWR VGND _05558_ _02550_ keymem.key_mem\[9\]\[21\] _05559_ sky130_fd_sc_hd__mux2_2
XFILLER_0_60_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22007_ VGND VPWR _06484_ _06405_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20199_ VGND VPWR _00874_ _05520_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_200_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1090 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_48_Left_316 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14760_ _09059_ _10226_ _09105_ _09046_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_23958_ VGND VPWR VPWR VGND clk _00451_ reset_n keymem.key_mem\[13\]\[79\] sky130_fd_sc_hd__dfrtp_2
X_11972_ VGND VPWR VGND VPWR _07542_ keymem.key_mem\[8\]\[0\] _07553_ _07570_ _07575_
+ _07574_ sky130_fd_sc_hd__a2111o_2
X_13711_ VGND VPWR VPWR VGND _09176_ _09182_ _09170_ _09183_ sky130_fd_sc_hd__or3_2
X_22909_ VGND VPWR VGND VPWR _06911_ _11457_ _03860_ _06884_ _11545_ sky130_fd_sc_hd__a211o_2
XFILLER_0_170_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14691_ VPWR VGND VGND VPWR _09127_ _10158_ _09211_ sky130_fd_sc_hd__nor2_2
XFILLER_0_196_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Right_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23889_ VGND VPWR VPWR VGND clk _00382_ reset_n keymem.key_mem\[13\]\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_211_461 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16430_ VPWR VGND VPWR VGND _02590_ _02592_ _02588_ _02589_ sky130_fd_sc_hd__or3b_2
XFILLER_0_131_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13642_ VGND VPWR _09114_ _09079_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25628_ VGND VPWR VPWR VGND clk _02121_ reset_n keymem.key_mem\[0\]\[85\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_170_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_168_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16361_ VPWR VGND VGND VPWR _11399_ _02524_ _11267_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_588 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13573_ VGND VPWR _09045_ _09034_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_211_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25559_ VGND VPWR VPWR VGND clk _02052_ reset_n keymem.key_mem\[0\]\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26_216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18100_ VPWR VGND VPWR VGND _04019_ _03970_ _09982_ sky130_fd_sc_hd__or2_2
X_15312_ VPWR VGND VGND VPWR _10773_ _10774_ _10770_ sky130_fd_sc_hd__nor2_2
X_12524_ VGND VPWR _08090_ _07761_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19080_ VGND VPWR VGND VPWR _04893_ keymem.key_mem_we _10836_ _04878_ _00382_ sky130_fd_sc_hd__a31o_2
XFILLER_0_13_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16292_ VPWR VGND VPWR VGND _02359_ _11518_ _02456_ _11476_ _02455_ sky130_fd_sc_hd__or4b_2
XPHY_EDGE_ROW_57_Left_325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_87_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18031_ VGND VPWR _03953_ _03952_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_81_366 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_240_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15243_ VGND VPWR VGND VPWR _10572_ _10569_ _10604_ _10478_ _10580_ _10706_ sky130_fd_sc_hd__o32a_2
X_12455_ VGND VPWR _08027_ _07534_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_81_388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15174_ VPWR VGND VGND VPWR _10575_ _10638_ _10478_ sky130_fd_sc_hd__nor2_2
X_12386_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[25\] _07963_ keymem.key_mem\[12\]\[25\]
+ _07788_ _07964_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_28_Right_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14125_ VGND VPWR VPWR VGND _09425_ _09443_ _09247_ _09596_ sky130_fd_sc_hd__or3_2
XFILLER_0_22_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19982_ VGND VPWR VPWR VGND _05400_ _11149_ keymem.key_mem\[10\]\[15\] _05407_ sky130_fd_sc_hd__mux2_2
XFILLER_0_10_639 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18933_ VPWR VGND _04770_ enc_block.block_w2_reg\[27\] enc_block.block_w3_reg\[23\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_14056_ VPWR VGND VPWR VGND _09528_ keymem.prev_key1_reg\[64\] sky130_fd_sc_hd__inv_2
XFILLER_0_219_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_24_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_103_1_Left_370 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_253_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13007_ VGND VPWR VGND VPWR _07584_ keymem.key_mem\[14\]\[84\] _08523_ _08525_ _08526_
+ _08480_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_94_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18864_ VPWR VGND VPWR VGND _04708_ _04664_ _04707_ enc_block.block_w2_reg\[11\]
+ _04602_ _00351_ sky130_fd_sc_hd__a221o_2
XFILLER_0_118_23 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_98_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17815_ VGND VPWR _00205_ _03805_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18795_ VPWR VGND _04646_ enc_block.block_w2_reg\[29\] enc_block.block_w3_reg\[21\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_234_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17746_ VGND VPWR VPWR VGND _03723_ _03761_ keymem.prev_key0_reg\[39\] _03762_ sky130_fd_sc_hd__mux2_2
X_14958_ VGND VPWR VGND VPWR enc_block.block_w2_reg\[13\] _09269_ _09021_ _10420_
+ _10422_ _10421_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_168_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Right_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_76_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13909_ VGND VPWR _09381_ _09380_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17677_ VGND VPWR _00158_ _03714_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_203_962 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14889_ VGND VPWR VGND VPWR _09173_ _09222_ _09113_ _09082_ _10354_ sky130_fd_sc_hd__o22a_2
X_19416_ VGND VPWR _00507_ _05104_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16628_ VPWR VGND VPWR VGND _02784_ key[156] _10286_ sky130_fd_sc_hd__or2_2
XFILLER_0_9_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_159_376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_1171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_174_335 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19347_ VGND VPWR VPWR VGND _05046_ _05058_ keymem.key_mem\[13\]\[112\] _05059_ sky130_fd_sc_hd__mux2_2
X_16559_ VPWR VGND VGND VPWR _02717_ _02718_ keylen sky130_fd_sc_hd__nor2_2
XFILLER_0_2_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_739 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_31_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19278_ VGND VPWR VPWR VGND _04993_ _05013_ keymem.key_mem\[13\]\[88\] _05014_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_249 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_154_1_Right_755 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_127_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_127_284 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_150_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18229_ VGND VPWR VGND VPWR _04136_ _03992_ _04133_ _04134_ _00288_ sky130_fd_sc_hd__a31o_2
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_644 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_142_243 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21240_ VGND VPWR VPWR VGND _06065_ _03443_ keymem.key_mem\[6\]\[93\] _06075_ sky130_fd_sc_hd__mux2_2
XFILLER_0_241_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_263 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21171_ VGND VPWR VPWR VGND _06029_ _03149_ keymem.key_mem\[6\]\[60\] _06039_ sky130_fd_sc_hd__mux2_2
XFILLER_0_159_74 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20122_ VGND VPWR VPWR VGND _05469_ _03347_ keymem.key_mem\[10\]\[82\] _05480_ sky130_fd_sc_hd__mux2_2
XFILLER_0_256_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_229_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20053_ VGND VPWR VPWR VGND _05435_ _03046_ keymem.key_mem\[10\]\[49\] _05444_ sky130_fd_sc_hd__mux2_2
XFILLER_0_238_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24930_ VGND VPWR VPWR VGND clk _01423_ reset_n keymem.key_mem\[5\]\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_209_Left_476 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24861_ VGND VPWR VPWR VGND clk _01354_ reset_n keymem.key_mem\[6\]\[86\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_704 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_55_Right_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23812_ VGND VPWR VPWR VGND clk _00305_ reset_n enc_block.block_w0_reg\[31\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_169_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24792_ VGND VPWR VPWR VGND clk _01285_ reset_n keymem.key_mem\[6\]\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_197_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23743_ keymem.prev_key0_reg\[99\] clk _00240_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_36_1033 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_67_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20955_ VGND VPWR _01226_ _05924_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_230_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_246_Right_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_221_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_221_792 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_113_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23674_ keymem.prev_key0_reg\[30\] clk _00171_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_48_330 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20886_ VPWR VGND keymem.key_mem\[7\]\[54\] _05888_ _05886_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_152_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25413_ VGND VPWR VPWR VGND clk _01906_ reset_n keymem.key_mem\[2\]\[126\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_179_1_Left_446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22625_ VGND VPWR _02038_ _06782_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_113_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_182 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_218_Left_485 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_147_2_Left_618 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25344_ VGND VPWR VPWR VGND clk _01837_ reset_n keymem.key_mem\[2\]\[57\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22556_ VGND VPWR _01988_ _06763_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_148_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1042 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_64_Right_64 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_84_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21507_ VGND VPWR _01486_ _06216_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25275_ VGND VPWR VPWR VGND clk _01768_ reset_n keymem.key_mem\[3\]\[116\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_1086 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_133_243 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22487_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[39\] _06707_ _06706_ _04933_ _01947_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_32_731 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24226_ VGND VPWR VPWR VGND clk _00719_ reset_n keymem.key_mem\[11\]\[91\] sky130_fd_sc_hd__dfrtp_2
X_12240_ VGND VPWR VGND VPWR _07830_ _07622_ keymem.key_mem\[13\]\[13\] _07827_ _07829_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_16_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1140 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21438_ VGND VPWR _01453_ _06180_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_210_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12171_ VGND VPWR enc_block.round_key\[8\] _07765_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21369_ VGND VPWR _01420_ _06144_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24157_ VGND VPWR VPWR VGND clk _00650_ reset_n keymem.key_mem\[11\]\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_47_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23108_ VGND VPWR _07032_ _06880_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24088_ VGND VPWR VPWR VGND clk _00581_ reset_n keymem.key_mem\[12\]\[81\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_120_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15930_ VGND VPWR _11386_ _11385_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_60_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_227_Left_494 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_159_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_66 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23039_ VGND VPWR _03224_ keylen _06990_ _03220_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_95_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_159_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15861_ VPWR VGND VPWR VGND _11192_ _11229_ _11207_ _11187_ _11317_ sky130_fd_sc_hd__or4_2
XFILLER_0_95_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17600_ VGND VPWR VGND VPWR _02829_ _02828_ _03658_ _10967_ sky130_fd_sc_hd__a21oi_2
X_14812_ VGND VPWR _10278_ _09523_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18580_ VGND VPWR _04453_ enc_block.block_w0_reg\[6\] _04452_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15792_ VGND VPWR VGND VPWR _11248_ _11215_ _11214_ keymem.prev_key1_reg\[16\] _08989_
+ _08983_ sky130_fd_sc_hd__a32o_2
XFILLER_0_118_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17531_ VGND VPWR VPWR VGND _09927_ _03597_ key[245] _03598_ sky130_fd_sc_hd__mux2_2
XFILLER_0_8_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14743_ _10207_ _10209_ _10206_ _10208_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_59_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11955_ VGND VPWR _07558_ _07557_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_93_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17462_ VGND VPWR VPWR VGND _03534_ keymem.key_mem\[14\]\[107\] _03538_ _03539_ sky130_fd_sc_hd__mux2_2
X_14674_ VPWR VGND VGND VPWR _10141_ _10108_ _10140_ sky130_fd_sc_hd__nand2_2
X_11886_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[14\] dec_new_block\[110\]
+ _07507_ sky130_fd_sc_hd__mux2_2
XFILLER_0_131_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16413_ VGND VPWR VGND VPWR _02574_ _11477_ _11340_ _11407_ _02575_ sky130_fd_sc_hd__a31o_2
X_19201_ VPWR VGND keymem.key_mem\[13\]\[58\] _04967_ _04961_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13625_ VGND VPWR _09097_ _09096_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_156_335 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_71_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17393_ VGND VPWR VGND VPWR _03478_ _02889_ _03477_ keylen _03479_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_131_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19132_ VGND VPWR VPWR VGND _04877_ _04922_ keymem.key_mem\[13\]\[33\] _04923_ sky130_fd_sc_hd__mux2_2
X_16344_ VGND VPWR VGND VPWR _02507_ _11365_ _11409_ _11427_ _11434_ _11222_ sky130_fd_sc_hd__a32o_2
XFILLER_0_109_251 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_183_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13556_ VPWR VGND VPWR VGND _08963_ _09027_ _08970_ _08957_ _09028_ sky130_fd_sc_hd__or4_2
XFILLER_0_32_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_878 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_89_16 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_54_377 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_67_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_124_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12507_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[35\] _07893_ _08074_ _08070_ _08075_
+ sky130_fd_sc_hd__o22a_2
X_19063_ VPWR VGND keymem.key_mem\[13\]\[3\] _04884_ _04880_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16275_ VGND VPWR VGND VPWR _02439_ _02436_ _11408_ _02437_ _02438_ sky130_fd_sc_hd__a211o_2
X_13487_ VPWR VGND VGND VPWR enc_block.block_w1_reg\[3\] enc_block.sword_ctr_reg\[0\]
+ _08959_ sky130_fd_sc_hd__or2b_2
X_18014_ VPWR VGND enc_block.round\[0\] _03941_ _07374_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_246_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15226_ VPWR VGND VGND VPWR _10449_ _10459_ _10689_ _10546_ _10539_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_124_265 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12438_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[29\] _07578_ keymem.key_mem\[8\]\[29\]
+ _07540_ _08012_ sky130_fd_sc_hd__a22o_2
XFILLER_0_65_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15157_ VGND VPWR _10620_ _10538_ _10621_ _10618_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_2_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12369_ VGND VPWR VGND VPWR _07949_ _07761_ keymem.key_mem\[11\]\[23\] _07948_ _07572_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_11_948 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_103_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14108_ VPWR VGND VGND VPWR _09563_ _09579_ _09380_ sky130_fd_sc_hd__nor2_2
XFILLER_0_107_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_193_2_Left_664 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_142_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15088_ VPWR VGND VGND VPWR _10493_ _10533_ _10551_ _10552_ sky130_fd_sc_hd__nor3_2
X_19965_ VGND VPWR _00763_ _05397_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_103_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18916_ VPWR VGND _04755_ enc_block.block_w0_reg\[9\] enc_block.block_w1_reg\[1\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_38_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14039_ VGND VPWR _09511_ _09510_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19896_ VGND VPWR _00732_ _05359_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_101_1160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18847_ VPWR VGND VGND VPWR _04693_ enc_block.block_w1_reg\[1\] enc_block.block_w1_reg\[2\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_253_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_257_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_175_1250 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_145_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_253_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18778_ VPWR VGND VPWR VGND block[35] _03979_ enc_block.block_w1_reg\[3\] _04138_
+ _04631_ sky130_fd_sc_hd__a22o_2
XFILLER_0_54_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17729_ VPWR VGND VPWR VGND _02859_ _03752_ keymem.prev_key0_reg\[31\] _03730_ _00172_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_49_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20740_ VGND VPWR VPWR VGND _05805_ _03600_ keymem.key_mem\[8\]\[117\] _05807_ sky130_fd_sc_hd__mux2_2
XFILLER_0_114_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20671_ VGND VPWR _01096_ _05770_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_45_300 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22410_ VGND VPWR _01908_ _06697_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_11_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23390_ VGND VPWR VGND VPWR _07262_ _04149_ _07095_ _07263_ enc_block.block_w3_reg\[18\]
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_247_1229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_184_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_942 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22341_ VGND VPWR VPWR VGND _06658_ _03466_ keymem.key_mem\[2\]\[96\] _06661_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_155_1_Right_756 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_225_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_264_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_474 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22272_ VGND VPWR VPWR VGND _06622_ _03183_ keymem.key_mem\[2\]\[63\] _06625_ sky130_fd_sc_hd__mux2_2
X_25060_ VGND VPWR VPWR VGND clk _01553_ reset_n keymem.key_mem\[4\]\[29\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_260_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21223_ VGND VPWR _01352_ _06066_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24011_ VGND VPWR VPWR VGND clk _00504_ reset_n keymem.key_mem\[12\]\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_121_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21154_ VGND VPWR _01319_ _06030_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_160_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20105_ VGND VPWR _00829_ _05471_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_10_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21085_ VGND VPWR VPWR VGND _05983_ _02409_ keymem.key_mem\[6\]\[19\] _05994_ sky130_fd_sc_hd__mux2_2
XFILLER_0_244_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_258_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20036_ VGND VPWR _05435_ _05388_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24913_ VGND VPWR VPWR VGND clk _01406_ reset_n keymem.key_mem\[5\]\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1166 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24844_ VGND VPWR VPWR VGND clk _01337_ reset_n keymem.key_mem\[6\]\[69\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_1199 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_232_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24775_ VGND VPWR VPWR VGND clk _01268_ reset_n keymem.key_mem\[6\]\[0\] sky130_fd_sc_hd__dfrtp_2
X_21987_ VGND VPWR VGND VPWR _06473_ keymem.key_mem_we _03119_ _06446_ _01709_ sky130_fd_sc_hd__a31o_2
X_23726_ keymem.prev_key0_reg\[82\] clk _00223_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_11740_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[5\] dec_new_block\[37\]
+ _07434_ sky130_fd_sc_hd__mux2_2
X_20938_ VGND VPWR _01218_ _05915_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_205_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11671_ VGND VPWR result[2] _07399_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23657_ keymem.prev_key0_reg\[13\] clk _00154_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20869_ VGND VPWR _01186_ _05878_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13410_ VPWR VGND VPWR VGND _08888_ keymem.key_mem\[3\]\[124\] _07844_ keymem.key_mem\[4\]\[124\]
+ _07914_ _08889_ sky130_fd_sc_hd__a221o_2
XFILLER_0_265_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22608_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[118\] _06777_ _06776_ _05071_ _02026_
+ sky130_fd_sc_hd__a22o_2
X_14390_ VGND VPWR VPWR VGND _09796_ key[2] _09860_ _09859_ _09857_ sky130_fd_sc_hd__o211a_2
X_23588_ VGND VPWR VPWR VGND clk _00089_ reset_n keymem.key_mem\[14\]\[77\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_889 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_349 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_51_303 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25327_ VGND VPWR VPWR VGND clk _01820_ reset_n keymem.key_mem\[2\]\[40\] sky130_fd_sc_hd__dfrtp_2
X_13341_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[117\] _07694_ keymem.key_mem\[10\]\[117\]
+ _07742_ _08827_ sky130_fd_sc_hd__a22o_2
XFILLER_0_64_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22539_ VGND VPWR VPWR VGND _06750_ keymem.key_mem\[1\]\[69\] _03235_ _06758_ sky130_fd_sc_hd__mux2_2
XFILLER_0_49_1246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16060_ VPWR VGND VGND VPWR _11514_ _11513_ _11395_ _11340_ _11357_ _11515_ sky130_fd_sc_hd__a311o_2
XFILLER_0_106_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25258_ VGND VPWR VPWR VGND clk _01751_ reset_n keymem.key_mem\[3\]\[99\] sky130_fd_sc_hd__dfrtp_2
X_13272_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[110\] _07842_ keymem.key_mem\[8\]\[110\]
+ _07542_ _08765_ sky130_fd_sc_hd__a22o_2
X_15011_ VPWR VGND VGND VPWR _10475_ _10440_ _10464_ sky130_fd_sc_hd__nand2_2
XFILLER_0_161_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24209_ VGND VPWR VPWR VGND clk _00702_ reset_n keymem.key_mem\[11\]\[74\] sky130_fd_sc_hd__dfrtp_2
X_12223_ VPWR VGND VPWR VGND _07813_ keymem.key_mem\[5\]\[12\] _07811_ keymem.key_mem\[8\]\[12\]
+ _07655_ _07814_ sky130_fd_sc_hd__a221o_2
XFILLER_0_267_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1340 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25189_ VGND VPWR VPWR VGND clk _01682_ reset_n keymem.key_mem\[3\]\[30\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_235_Left_502 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12154_ VGND VPWR VGND VPWR _07737_ keymem.key_mem\[1\]\[7\] _07741_ _07747_ _07750_
+ _07749_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_236_604 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_124_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19750_ VGND VPWR _00662_ _05283_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16962_ VGND VPWR VPWR VGND _03084_ keymem.key_mem\[14\]\[54\] _03091_ _03092_ sky130_fd_sc_hd__mux2_2
X_12085_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[4\] _07620_ keymem.key_mem\[8\]\[4\]
+ _07654_ _07684_ sky130_fd_sc_hd__a22o_2
XFILLER_0_159_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18701_ VGND VPWR _04561_ enc_block.block_w2_reg\[20\] enc_block.block_w0_reg\[4\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15913_ VPWR VGND VPWR VGND _11192_ _11202_ _11197_ _11225_ _11369_ sky130_fd_sc_hd__or4_2
XFILLER_0_95_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16893_ VGND VPWR _03029_ _09987_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19681_ VGND VPWR _05247_ _05246_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_246_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1100 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15844_ VGND VPWR VGND VPWR _11300_ _11299_ _11285_ _11277_ sky130_fd_sc_hd__and3b_2
X_18632_ VPWR VGND VGND VPWR _04499_ _04500_ _04478_ sky130_fd_sc_hd__nor2_2
XFILLER_0_95_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_692 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_246_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_188_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15775_ _11224_ _11231_ _11222_ _11230_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_18563_ VPWR VGND VPWR VGND _04438_ _04434_ _04436_ sky130_fd_sc_hd__or2_2
X_12987_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[82\] _07613_ keymem.key_mem\[10\]\[82\]
+ _08193_ _08508_ sky130_fd_sc_hd__a22o_2
XFILLER_0_8_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_244_Left_511 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_262_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17514_ VGND VPWR VPWR VGND _10378_ _02402_ key[243] _03583_ sky130_fd_sc_hd__mux2_2
X_14726_ VPWR VGND VPWR VGND _10192_ _09638_ _10145_ key[133] _09544_ _10193_ sky130_fd_sc_hd__a221o_2
X_18494_ VPWR VGND VPWR VGND _04376_ _04372_ _04374_ sky130_fd_sc_hd__or2_2
X_11938_ VGND VPWR _07541_ _07540_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_262_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17445_ VPWR VGND _09533_ _03524_ _03523_ VPWR VGND sky130_fd_sc_hd__and2_2
X_14657_ VGND VPWR VGND VPWR _09388_ _09355_ _09312_ _09408_ _10124_ sky130_fd_sc_hd__o22a_2
XFILLER_0_156_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11869_ VGND VPWR result[101] _07498_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_717 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_6_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13608_ VGND VPWR _09080_ _09079_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17376_ VPWR VGND key[224] _03464_ _09868_ VPWR VGND sky130_fd_sc_hd__and2_2
X_14588_ VGND VPWR VGND VPWR _10040_ _10055_ _10056_ _10033_ _10046_ sky130_fd_sc_hd__nor4_2
XFILLER_0_171_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16327_ VPWR VGND VPWR VGND keymem.prev_key1_reg\[53\] _02490_ _02488_ _02489_ sky130_fd_sc_hd__or3b_2
X_19115_ VPWR VGND keymem.key_mem\[13\]\[26\] _04913_ _04903_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13539_ VPWR VGND VGND VPWR _09011_ _09009_ _09010_ sky130_fd_sc_hd__nand2_2
XFILLER_0_40_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_539 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_67_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19046_ VPWR VGND VPWR VGND _04870_ _04505_ enc_block.block_w2_reg\[31\] _04504_
+ _04871_ sky130_fd_sc_hd__a22o_2
X_16258_ VGND VPWR VGND VPWR _11219_ _11375_ _11379_ _11320_ _02422_ sky130_fd_sc_hd__o22a_2
XFILLER_0_42_358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_67_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15209_ VGND VPWR _10672_ _10439_ _10483_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_253_Left_520 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_258_217 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_207_1257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16189_ VGND VPWR VGND VPWR _11283_ _11469_ _11395_ _02353_ _02354_ sky130_fd_sc_hd__o22a_2
XFILLER_0_3_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_380 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_239_442 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19948_ VGND VPWR _05388_ _05387_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_208_851 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_78_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19879_ VGND VPWR VPWR VGND _05350_ keymem.key_mem\[11\]\[96\] _03466_ _05351_ sky130_fd_sc_hd__mux2_2
XFILLER_0_65_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_177_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21910_ VGND VPWR _06432_ _06403_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_78_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22890_ VGND VPWR VPWR VGND _06878_ _10745_ keymem.prev_key1_reg\[9\] _06900_ sky130_fd_sc_hd__mux2_2
XFILLER_0_74_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_662 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21841_ VGND VPWR VPWR VGND _06388_ _03620_ keymem.key_mem\[4\]\[120\] _06393_ sky130_fd_sc_hd__mux2_2
XFILLER_0_172_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24560_ VGND VPWR VPWR VGND clk _01053_ reset_n keymem.key_mem\[8\]\[41\] sky130_fd_sc_hd__dfrtp_2
X_21772_ VGND VPWR VPWR VGND _06355_ _03392_ keymem.key_mem\[4\]\[87\] _06357_ sky130_fd_sc_hd__mux2_2
XFILLER_0_210_559 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_114_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23511_ VGND VPWR VPWR VGND clk _00012_ reset_n keymem.key_mem\[14\]\[0\] sky130_fd_sc_hd__dfrtp_2
X_20723_ VGND VPWR VPWR VGND _05794_ _03550_ keymem.key_mem\[8\]\[109\] _05798_ sky130_fd_sc_hd__mux2_2
X_24491_ VGND VPWR VPWR VGND clk _00984_ reset_n keymem.key_mem\[9\]\[100\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_11_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23442_ VGND VPWR VGND VPWR _03959_ block[24] _07309_ _07308_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_149_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20654_ VGND VPWR VPWR VGND _05761_ _03295_ keymem.key_mem\[8\]\[76\] _05762_ sky130_fd_sc_hd__mux2_2
XFILLER_0_188_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_11_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_303 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23373_ VGND VPWR _07247_ enc_block.block_w2_reg\[1\] _07246_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20585_ VGND VPWR VPWR VGND _05725_ _02985_ keymem.key_mem\[8\]\[43\] _05726_ sky130_fd_sc_hd__mux2_2
XFILLER_0_85_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25112_ VGND VPWR VPWR VGND clk _01605_ reset_n keymem.key_mem\[4\]\[81\] sky130_fd_sc_hd__dfrtp_2
X_22324_ VGND VPWR VPWR VGND _06647_ _03401_ keymem.key_mem\[2\]\[88\] _06652_ sky130_fd_sc_hd__mux2_2
XFILLER_0_103_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_156_1_Right_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_85_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25043_ VGND VPWR VPWR VGND clk _01536_ reset_n keymem.key_mem\[4\]\[12\] sky130_fd_sc_hd__dfrtp_2
X_22255_ VGND VPWR VPWR VGND _06611_ _03099_ keymem.key_mem\[2\]\[55\] _06616_ sky130_fd_sc_hd__mux2_2
X_21206_ VGND VPWR _01344_ _06057_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22186_ VGND VPWR VPWR VGND _06578_ _02607_ keymem.key_mem\[2\]\[22\] _06580_ sky130_fd_sc_hd__mux2_2
XFILLER_0_121_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_946 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21137_ VGND VPWR _01311_ _06021_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_199_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_22_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21068_ VGND VPWR VGND VPWR keymem.round_ctr_reg\[3\] keymem.round_ctr_reg\[2\] _05385_
+ _05985_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_96_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_156_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1008 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_233_629 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_254_990 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20019_ VGND VPWR _00788_ _05426_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12910_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[74\] _08259_ _08438_ _08434_ _08439_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_260_437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13890_ VGND VPWR _09362_ _09317_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_96_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_21_Left_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_57_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24827_ VGND VPWR VPWR VGND clk _01320_ reset_n keymem.key_mem\[6\]\[52\] sky130_fd_sc_hd__dfrtp_2
X_12841_ VGND VPWR enc_block.round_key\[67\] _08376_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_214_887 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_236_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15560_ VGND VPWR VPWR VGND _10993_ _11018_ _07386_ _11019_ sky130_fd_sc_hd__or3_2
X_12772_ VGND VPWR enc_block.round_key\[60\] _08314_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24758_ VGND VPWR VPWR VGND clk _01251_ reset_n keymem.key_mem\[7\]\[111\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_56_406 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14511_ VPWR VGND VGND VPWR _09973_ _09975_ _09977_ _09979_ _09980_ sky130_fd_sc_hd__and4b_2
X_11723_ VGND VPWR result[28] _07425_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23709_ keymem.prev_key0_reg\[65\] clk _00206_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_132_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15491_ VGND VPWR VGND VPWR _10482_ _10668_ _10629_ _10527_ _10951_ sky130_fd_sc_hd__o22a_2
X_24689_ VGND VPWR VPWR VGND clk _01182_ reset_n keymem.key_mem\[7\]\[42\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17230_ _11535_ _03333_ _03332_ _11536_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_14442_ VPWR VGND VGND VPWR _09381_ _09911_ _09268_ sky130_fd_sc_hd__nor2_2
XFILLER_0_167_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_37_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11654_ VGND VPWR VGND VPWR _07390_ _07389_ _00002_ keymem.round_ctr_rst sky130_fd_sc_hd__o21a_2
XFILLER_0_153_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17161_ VGND VPWR VGND VPWR _10818_ _10817_ _03271_ keymem.prev_key0_reg\[74\] sky130_fd_sc_hd__a21oi_2
X_14373_ VGND VPWR VGND VPWR _09029_ _09050_ _09684_ _09082_ _09843_ sky130_fd_sc_hd__o22a_2
XFILLER_0_49_1021 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_24_325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_30_Left_298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16112_ VPWR VGND VGND VPWR _11367_ _11566_ _11239_ sky130_fd_sc_hd__nor2_2
XFILLER_0_52_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13324_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[115\] _08714_ _08811_ _08807_ _08812_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_101_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_243_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17092_ VGND VPWR VPWR VGND _03185_ keymem.key_mem\[14\]\[66\] _03209_ _03210_ sky130_fd_sc_hd__mux2_2
XFILLER_0_208_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16043_ VGND VPWR VGND VPWR _11460_ _11497_ _11498_ _11252_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_33_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13255_ VGND VPWR VGND VPWR _08750_ _07839_ keymem.key_mem\[11\]\[108\] _08747_ _08749_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_161_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12206_ VGND VPWR VGND VPWR _07753_ keymem.key_mem\[8\]\[11\] _07795_ _07797_ _07798_
+ _07616_ sky130_fd_sc_hd__a2111o_2
X_13186_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[102\] _08016_ keymem.key_mem\[6\]\[102\]
+ _07908_ _08687_ sky130_fd_sc_hd__a22o_2
XFILLER_0_20_564 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_104_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19802_ VGND VPWR _00687_ _05310_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_237_946 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12137_ VGND VPWR _07733_ _07732_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_104_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17994_ VGND VPWR VGND VPWR _03928_ _03927_ _03675_ _03625_ sky130_fd_sc_hd__and3b_2
XFILLER_0_40_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19733_ VGND VPWR _00654_ _05274_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12068_ VGND VPWR _07668_ _07667_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16945_ VGND VPWR _00064_ _03076_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_223_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_174_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19664_ VGND VPWR VPWR VGND _05227_ _05083_ keymem.key_mem\[12\]\[124\] _05236_ sky130_fd_sc_hd__mux2_2
X_16876_ VPWR VGND VGND VPWR _03014_ key[174] _02875_ sky130_fd_sc_hd__nand2_2
XFILLER_0_216_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_254_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18615_ VPWR VGND _04485_ _04484_ enc_block.round_key\[82\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_260_971 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15827_ VGND VPWR _11283_ _11282_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19595_ VPWR VGND keymem.key_mem\[12\]\[91\] _05200_ _05094_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_215_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_59_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15758_ VGND VPWR VGND VPWR enc_block.block_w1_reg\[16\] _08985_ _10387_ _11212_
+ _11214_ _11213_ sky130_fd_sc_hd__a2111o_2
X_18546_ VPWR VGND VGND VPWR _04380_ _04423_ _04107_ sky130_fd_sc_hd__nor2_2
XFILLER_0_248_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14709_ VPWR VGND VGND VPWR _09127_ _10176_ _09222_ sky130_fd_sc_hd__nor2_2
X_18477_ VPWR VGND _04361_ _04360_ enc_block.round_key\[68\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15689_ VGND VPWR VPWR VGND _11146_ _09717_ _11111_ _11144_ _09721_ sky130_fd_sc_hd__o31a_2
XFILLER_0_74_236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17428_ VGND VPWR VGND VPWR _03508_ _02943_ _03509_ keylen sky130_fd_sc_hd__a21oi_2
XFILLER_0_117_349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17359_ VGND VPWR VGND VPWR key[94] _08937_ _03448_ _03447_ _03449_ sky130_fd_sc_hd__o22a_2
XFILLER_0_16_859 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_43_656 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20370_ VGND VPWR VPWR VGND _05602_ _03245_ keymem.key_mem\[9\]\[70\] _05612_ sky130_fd_sc_hd__mux2_2
XFILLER_0_261_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_63_1018 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19029_ VGND VPWR _04856_ _04647_ _04855_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22040_ VPWR VGND keymem.key_mem\[3\]\[82\] _06502_ _06484_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_140_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_80_1_Right_681 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_55_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_188_1_Left_455 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23991_ VGND VPWR VPWR VGND clk _00484_ reset_n keymem.key_mem\[13\]\[112\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_214_117 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_199_319 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_156_2_Left_627 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25730_ keymem.prev_key1_reg\[46\] clk _02223_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_39_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22942_ VGND VPWR VGND VPWR _06933_ _02775_ _06891_ _02785_ _06892_ sky130_fd_sc_hd__a211o_2
XFILLER_0_78_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_40 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25661_ VGND VPWR VPWR VGND clk _02154_ reset_n keymem.key_mem\[0\]\[118\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_92_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22873_ VPWR VGND VGND VPWR _06881_ _06889_ keymem.prev_key1_reg\[3\] sky130_fd_sc_hd__nor2_2
XFILLER_0_218_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24612_ VGND VPWR VPWR VGND clk _01105_ reset_n keymem.key_mem\[8\]\[93\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_210_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21824_ VGND VPWR VPWR VGND _06377_ _03567_ keymem.key_mem\[4\]\[112\] _06384_ sky130_fd_sc_hd__mux2_2
X_25592_ VGND VPWR VPWR VGND clk _02085_ reset_n keymem.key_mem\[0\]\[49\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_167_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_151_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24543_ VGND VPWR VPWR VGND clk _01036_ reset_n keymem.key_mem\[8\]\[24\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_65_214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21755_ VGND VPWR VPWR VGND _06344_ _03321_ keymem.key_mem\[4\]\[79\] _06348_ sky130_fd_sc_hd__mux2_2
XFILLER_0_108_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20706_ VGND VPWR VPWR VGND _05783_ _03499_ keymem.key_mem\[8\]\[101\] _05789_ sky130_fd_sc_hd__mux2_2
XFILLER_0_135_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24474_ VGND VPWR VPWR VGND clk _00967_ reset_n keymem.key_mem\[9\]\[83\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_135_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21686_ VGND VPWR VPWR VGND _06308_ _03015_ keymem.key_mem\[4\]\[46\] _06312_ sky130_fd_sc_hd__mux2_2
XFILLER_0_149_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_686 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23425_ VGND VPWR VGND VPWR _03958_ block[22] _07293_ _07294_ sky130_fd_sc_hd__a21o_2
X_20637_ VPWR VGND VGND VPWR _05676_ _05753_ keymem.key_mem\[8\]\[68\] sky130_fd_sc_hd__nor2_2
XFILLER_0_18_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_149_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23356_ VGND VPWR _07232_ enc_block.block_w2_reg\[7\] _07231_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20568_ VGND VPWR VPWR VGND _05714_ _02903_ keymem.key_mem\[8\]\[35\] _05717_ sky130_fd_sc_hd__mux2_2
XFILLER_0_264_1170 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_15_881 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22307_ VGND VPWR VPWR VGND _06634_ _03329_ keymem.key_mem\[2\]\[80\] _06643_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_157_1_Right_758 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23287_ VPWR VGND VGND VPWR _07170_ _07166_ _07168_ sky130_fd_sc_hd__nand2_2
X_20499_ VGND VPWR VPWR VGND _05680_ _09861_ keymem.key_mem\[8\]\[2\] _05681_ sky130_fd_sc_hd__mux2_2
XFILLER_0_260_1067 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13040_ VPWR VGND VPWR VGND _08555_ keymem.key_mem\[9\]\[87\] _07672_ keymem.key_mem\[8\]\[87\]
+ _08265_ _08556_ sky130_fd_sc_hd__a221o_2
X_25026_ VGND VPWR VPWR VGND clk _01519_ reset_n keymem.key_mem\[5\]\[123\] sky130_fd_sc_hd__dfrtp_2
X_22238_ VGND VPWR VPWR VGND _06600_ _03024_ keymem.key_mem\[2\]\[47\] _06607_ sky130_fd_sc_hd__mux2_2
XFILLER_0_162_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22169_ VGND VPWR VPWR VGND _06565_ _11098_ keymem.key_mem\[2\]\[14\] _06571_ sky130_fd_sc_hd__mux2_2
XFILLER_0_219_979 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_88_2_Left_559 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14991_ VGND VPWR _10455_ _10454_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_195_1264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13942_ _09412_ _09414_ _09406_ _09413_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_57_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16730_ VGND VPWR VGND VPWR _09634_ _09633_ _02880_ _02881_ sky130_fd_sc_hd__a21o_2
XFILLER_0_260_223 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_57_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16661_ VGND VPWR VGND VPWR keymem.rcon_logic.tmp_rcon\[7\] _02586_ _02572_ _02815_
+ sky130_fd_sc_hd__nand3b_2
X_13873_ VGND VPWR _09344_ _09327_ _09345_ _09330_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_202_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15612_ VPWR VGND VGND VPWR _10519_ _10536_ _10522_ _10667_ _11070_ _10491_ sky130_fd_sc_hd__o221a_2
X_18400_ VGND VPWR VGND VPWR _10261_ _10243_ _04073_ _04292_ sky130_fd_sc_hd__a21o_2
XFILLER_0_214_695 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_198_374 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12824_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[66\] _07845_ keymem.key_mem\[12\]\[66\]
+ _07788_ _08361_ sky130_fd_sc_hd__a22o_2
XFILLER_0_158_216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19380_ VPWR VGND keymem.key_mem_we _05081_ _03640_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16592_ VGND VPWR VGND VPWR _02748_ _10360_ _02746_ _02747_ _02749_ sky130_fd_sc_hd__a31o_2
XFILLER_0_232_1158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15543_ VGND VPWR VGND VPWR _10489_ _10411_ _11002_ _10507_ sky130_fd_sc_hd__a21oi_2
X_18331_ VPWR VGND VPWR VGND _04229_ block[119] _04213_ enc_block.block_w1_reg\[23\]
+ _04171_ _04230_ sky130_fd_sc_hd__a221o_2
X_12755_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[59\] _07818_ keymem.key_mem\[4\]\[59\]
+ _07854_ _08299_ sky130_fd_sc_hd__a22o_2
X_11706_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[20\] dec_new_block\[20\]
+ _07417_ sky130_fd_sc_hd__mux2_2
X_18262_ VPWR VGND VPWR VGND _04166_ block[113] _04076_ enc_block.block_w1_reg\[17\]
+ _04007_ _04167_ sky130_fd_sc_hd__a221o_2
X_15474_ VPWR VGND VPWR VGND _10710_ _10786_ _10933_ _10578_ _10934_ sky130_fd_sc_hd__or4_2
XFILLER_0_126_102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12686_ VPWR VGND VPWR VGND _08236_ keymem.key_mem\[11\]\[52\] _08011_ keymem.key_mem\[1\]\[52\]
+ _07671_ _08237_ sky130_fd_sc_hd__a221o_2
XFILLER_0_167_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14425_ VPWR VGND VGND VPWR _09565_ _09894_ _09353_ sky130_fd_sc_hd__nor2_2
XFILLER_0_25_612 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17213_ VPWR VGND VPWR VGND keymem.prev_key0_reg\[79\] _03318_ _11624_ _11144_ sky130_fd_sc_hd__or3b_2
XFILLER_0_126_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18193_ VGND VPWR VGND VPWR _04104_ _04103_ _04102_ _04101_ sky130_fd_sc_hd__and3b_2
X_11637_ VPWR VGND VGND VPWR _07376_ enc_block.sword_ctr_reg\[0\] enc_block.sword_ctr_reg\[1\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_25_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_4_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17144_ VGND VPWR _09513_ key[72] _03256_ _10366_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_14356_ VPWR VGND VPWR VGND _09824_ _09823_ _09825_ _09686_ _09826_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_68_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_107_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_188_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_486 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_97_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13307_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[114\] _07685_ keymem.key_mem\[4\]\[114\]
+ _07636_ _08796_ sky130_fd_sc_hd__a22o_2
XFILLER_0_12_328 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17075_ VGND VPWR VPWR VGND _03185_ keymem.key_mem\[14\]\[64\] _03194_ _03195_ sky130_fd_sc_hd__mux2_2
X_14287_ VGND VPWR VGND VPWR _09415_ _09404_ _09476_ _09756_ _09757_ sky130_fd_sc_hd__a31o_2
XFILLER_0_29_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16026_ VPWR VGND VPWR VGND _11478_ _11480_ _11479_ _11476_ _11481_ sky130_fd_sc_hd__or4_2
XFILLER_0_122_385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13238_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[107\] _07656_ keymem.key_mem\[11\]\[107\]
+ _07658_ _08734_ sky130_fd_sc_hd__a22o_2
XFILLER_0_20_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_423 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13169_ VPWR VGND VPWR VGND _08671_ keymem.key_mem\[14\]\[100\] _07666_ keymem.key_mem\[6\]\[100\]
+ _07818_ _08672_ sky130_fd_sc_hd__a221o_2
XFILLER_0_198_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1057 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_264_562 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_178_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17977_ VGND VPWR _00256_ _03916_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_174_1304 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_97_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19716_ VGND VPWR _00646_ _05265_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_139_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16928_ VPWR VGND VPWR VGND _03061_ _11624_ _03059_ _02396_ _03060_ _09721_ sky130_fd_sc_hd__o311a_2
XFILLER_0_252_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_119_1_Right_720 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_75_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19647_ VGND VPWR _05227_ _05091_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16859_ VGND VPWR VPWR VGND _02986_ keymem.key_mem\[14\]\[44\] _02998_ _02999_ sky130_fd_sc_hd__mux2_2
XFILLER_0_219_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1312 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19578_ VGND VPWR VGND VPWR _05191_ keymem.key_mem_we _03347_ _05187_ _00582_ sky130_fd_sc_hd__a31o_2
XFILLER_0_62_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18529_ VPWR VGND VPWR VGND _04407_ _04291_ _04406_ enc_block.block_w1_reg\[9\] _04317_
+ _00317_ sky130_fd_sc_hd__a221o_2
XFILLER_0_87_383 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_47_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_62_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21540_ VGND VPWR VPWR VGND _06231_ _03533_ keymem.key_mem\[5\]\[106\] _06234_ sky130_fd_sc_hd__mux2_2
XFILLER_0_117_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1110 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_63_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1143 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_69_1249 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21471_ VGND VPWR VPWR VGND _06196_ _03267_ keymem.key_mem\[5\]\[73\] _06198_ sky130_fd_sc_hd__mux2_2
X_23210_ VGND VPWR _07100_ _07098_ _07099_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_248_1176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20422_ VGND VPWR _00978_ _05639_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_86_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1029 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24190_ VGND VPWR VPWR VGND clk _00683_ reset_n keymem.key_mem\[11\]\[55\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_47_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_475 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_226_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23141_ VGND VPWR VGND VPWR _07052_ _03794_ _03537_ _07053_ sky130_fd_sc_hd__a21o_2
X_20353_ VGND VPWR _00945_ _05603_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_226_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23072_ VGND VPWR _07010_ _06881_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20284_ VGND VPWR VPWR VGND _05558_ _02812_ keymem.key_mem\[9\]\[29\] _05567_ sky130_fd_sc_hd__mux2_2
XFILLER_0_41_1102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_199_Right_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_1282 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22023_ VGND VPWR _01726_ _06492_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_81_1_Right_682 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_80_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_787 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_215_415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_259_1283 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_157_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23974_ VGND VPWR VPWR VGND clk _00467_ reset_n keymem.key_mem\[13\]\[95\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_199_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_118_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25713_ keymem.prev_key1_reg\[29\] clk _02206_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_39_1042 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22925_ VGND VPWR VGND VPWR _02649_ _02648_ _02659_ _06921_ sky130_fd_sc_hd__a21o_2
XFILLER_0_233_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25644_ VGND VPWR VPWR VGND clk _02137_ reset_n keymem.key_mem\[0\]\[101\] sky130_fd_sc_hd__dfrtp_2
X_22856_ VGND VPWR VGND VPWR _06876_ _05824_ _02175_ keymem.round_ctr_rst sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_155_1292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21807_ VGND VPWR VPWR VGND _06366_ _03518_ keymem.key_mem\[4\]\[104\] _06375_ sky130_fd_sc_hd__mux2_2
XFILLER_0_91_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25575_ VGND VPWR VPWR VGND clk _02068_ reset_n keymem.key_mem\[0\]\[32\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_78_394 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22787_ VGND VPWR _02128_ _06854_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_93_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12540_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[38\] _07893_ _08104_ _08098_ _08105_
+ sky130_fd_sc_hd__o22a_2
X_24526_ VGND VPWR VPWR VGND clk _01019_ reset_n keymem.key_mem\[8\]\[7\] sky130_fd_sc_hd__dfrtp_2
X_21738_ VGND VPWR VPWR VGND _06330_ _03251_ keymem.key_mem\[4\]\[71\] _06339_ sky130_fd_sc_hd__mux2_2
XFILLER_0_52_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_932 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24457_ VGND VPWR VPWR VGND clk _00950_ reset_n keymem.key_mem\[9\]\[66\] sky130_fd_sc_hd__dfrtp_2
X_12471_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[32\] _07600_ keymem.key_mem\[1\]\[32\]
+ _07799_ _08042_ sky130_fd_sc_hd__a22o_2
X_21669_ VGND VPWR VPWR VGND _06297_ _02934_ keymem.key_mem\[4\]\[38\] _06303_ sky130_fd_sc_hd__mux2_2
X_14210_ VGND VPWR VPWR VGND _09157_ _09033_ _09086_ _09681_ sky130_fd_sc_hd__or3_2
X_23408_ VPWR VGND VGND VPWR _07278_ _07279_ _04382_ sky130_fd_sc_hd__nor2_2
X_15190_ VGND VPWR VPWR VGND keymem.round_ctr_reg\[0\] _10653_ _09239_ _10654_ sky130_fd_sc_hd__mux2_2
XFILLER_0_34_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24388_ VGND VPWR VPWR VGND clk _00881_ reset_n keymem.key_mem\[10\]\[125\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_244_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14141_ VGND VPWR VGND VPWR _09416_ _09373_ _09495_ _09612_ sky130_fd_sc_hd__a21o_2
X_23339_ VGND VPWR VGND VPWR _07217_ _03955_ _07216_ _07215_ sky130_fd_sc_hd__o21a_2
XFILLER_0_205_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14072_ VGND VPWR _09543_ _08928_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_162_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_158_1_Right_759 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_205_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13023_ VGND VPWR enc_block.round_key\[85\] _08540_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25009_ VGND VPWR VPWR VGND clk _01502_ reset_n keymem.key_mem\[5\]\[106\] sky130_fd_sc_hd__dfrtp_2
X_17900_ VGND VPWR _03864_ _03679_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_63_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_197_1315 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18880_ VGND VPWR VGND VPWR _04723_ _04505_ _04722_ _04721_ sky130_fd_sc_hd__o21a_2
XFILLER_0_238_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17831_ VGND VPWR VPWR VGND _03814_ _03816_ keymem.prev_key0_reg\[69\] _03817_ sky130_fd_sc_hd__mux2_2
XFILLER_0_140_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_234_724 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_234_735 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17762_ VGND VPWR VPWR VGND _03763_ _03003_ keymem.prev_key0_reg\[45\] _03772_ sky130_fd_sc_hd__mux2_2
X_14974_ VGND VPWR VGND VPWR _10414_ _10411_ _10438_ _10437_ sky130_fd_sc_hd__a21oi_2
X_19501_ VPWR VGND keymem.key_mem\[12\]\[47\] _05150_ _05128_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16713_ VGND VPWR VPWR VGND _02864_ _09508_ _08931_ _02865_ sky130_fd_sc_hd__or3_2
X_13925_ VGND VPWR _09397_ _09322_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17693_ VGND VPWR VPWR VGND _03719_ key[151] keymem.prev_key1_reg\[23\] _03725_ sky130_fd_sc_hd__mux2_2
XFILLER_0_254_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19432_ VPWR VGND keymem.key_mem\[12\]\[15\] _05113_ _05102_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13856_ VGND VPWR _09328_ _09280_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16644_ VGND VPWR VGND VPWR _02536_ _11301_ _02799_ keymem.rcon_logic.tmp_rcon\[6\]
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_254_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12807_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[64\] _08050_ keymem.key_mem\[4\]\[64\]
+ _07841_ _08346_ sky130_fd_sc_hd__a22o_2
XFILLER_0_70_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_130_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19363_ VGND VPWR VPWR VGND _05067_ _05069_ keymem.key_mem\[13\]\[117\] _05070_ sky130_fd_sc_hd__mux2_2
XFILLER_0_29_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13787_ VPWR VGND VPWR VGND _09259_ enc_block.block_w0_reg\[26\] _08995_ sky130_fd_sc_hd__or2_2
XFILLER_0_134_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16575_ VGND VPWR VGND VPWR _02725_ _02724_ _02733_ keymem.prev_key1_reg\[122\] sky130_fd_sc_hd__a21oi_2
X_18314_ VGND VPWR _04214_ enc_block.block_w3_reg\[6\] enc_block.block_w1_reg\[21\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15526_ VGND VPWR VGND VPWR _10545_ _10573_ _10557_ _10587_ _10985_ sky130_fd_sc_hd__o22a_2
X_12738_ VPWR VGND VPWR VGND _08283_ keymem.key_mem\[14\]\[57\] _07685_ keymem.key_mem\[9\]\[57\]
+ _07716_ _08284_ sky130_fd_sc_hd__a221o_2
XFILLER_0_31_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19294_ VPWR VGND keymem.key_mem\[13\]\[95\] _05023_ _04879_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_139_293 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18245_ VGND VPWR _04151_ _03976_ _00289_ _04137_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_15457_ VPWR VGND VGND VPWR _10031_ _10917_ _10003_ sky130_fd_sc_hd__nor2_2
X_12669_ VGND VPWR enc_block.round_key\[50\] _08221_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14408_ VGND VPWR VGND VPWR _09876_ _09468_ _09360_ _09464_ _09877_ sky130_fd_sc_hd__a31o_2
XFILLER_0_113_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15388_ VPWR VGND VPWR VGND _10847_ _10848_ _10849_ _10438_ _10761_ sky130_fd_sc_hd__or4b_2
X_18176_ VPWR VGND _04088_ enc_block.block_w2_reg\[9\] enc_block.block_w3_reg\[1\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_52_261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_29_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14339_ VPWR VGND VGND VPWR _09083_ _09809_ _09136_ sky130_fd_sc_hd__nor2_2
X_17127_ VGND VPWR _03240_ _03238_ _03241_ _03239_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_204_1013 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_141_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_208_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17058_ _02854_ _03179_ _03178_ _02855_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_180_1385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16009_ VGND VPWR _11464_ _11302_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_81_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_141_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_265_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_209_275 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_57_96 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_768 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_252_565 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_174_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20971_ VGND VPWR _01234_ _05932_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_73_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_206_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22710_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[48\] _06820_ _06819_ _04950_ _02084_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_79_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23690_ keymem.prev_key0_reg\[46\] clk _00187_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_152_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_220_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22641_ VGND VPWR VPWR VGND _06785_ keymem.key_mem\[0\]\[9\] _10747_ _06792_ sky130_fd_sc_hd__mux2_2
XFILLER_0_152_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25360_ VGND VPWR VPWR VGND clk _01853_ reset_n keymem.key_mem\[2\]\[73\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_230_Right_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22572_ VGND VPWR _01998_ _06769_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_192_347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24311_ VGND VPWR VPWR VGND clk _00804_ reset_n keymem.key_mem\[10\]\[48\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_267_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21523_ VGND VPWR VPWR VGND _06220_ _03480_ keymem.key_mem\[5\]\[98\] _06225_ sky130_fd_sc_hd__mux2_2
X_25291_ VGND VPWR VPWR VGND clk _01784_ reset_n keymem.key_mem\[2\]\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_145_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24242_ VGND VPWR VPWR VGND clk _00735_ reset_n keymem.key_mem\[11\]\[107\] sky130_fd_sc_hd__dfrtp_2
X_21454_ VGND VPWR VPWR VGND _06184_ _03202_ keymem.key_mem\[5\]\[65\] _06189_ sky130_fd_sc_hd__mux2_2
XFILLER_0_146_1214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_263_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20405_ VGND VPWR _00970_ _05630_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24173_ VGND VPWR VPWR VGND clk _00666_ reset_n keymem.key_mem\[11\]\[38\] sky130_fd_sc_hd__dfrtp_2
X_21385_ VGND VPWR VPWR VGND _06151_ _02873_ keymem.key_mem\[5\]\[32\] _06153_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23124_ VGND VPWR VPWR VGND _07032_ _07041_ keymem.prev_key1_reg\[101\] _07042_ sky130_fd_sc_hd__mux2_2
X_20336_ VGND VPWR _00937_ _05594_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_163_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_222_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_990 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_12_692 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_60_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23055_ VPWR VGND VGND VPWR _06881_ _07000_ keymem.prev_key1_reg\[74\] sky130_fd_sc_hd__nor2_2
X_20267_ VGND VPWR _05558_ _05534_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_101_388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_82_1_Right_683 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22006_ VGND VPWR _01718_ _06483_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_228_562 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20198_ VGND VPWR VPWR VGND _05515_ _03607_ keymem.key_mem\[10\]\[118\] _05520_ sky130_fd_sc_hd__mux2_2
XFILLER_0_200_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_216_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11971_ VGND VPWR _07574_ _07573_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23957_ VGND VPWR VPWR VGND clk _00450_ reset_n keymem.key_mem\[13\]\[78\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13710_ VGND VPWR VGND VPWR _09182_ _09181_ _09180_ _09179_ sky130_fd_sc_hd__o21a_2
X_22908_ VGND VPWR _02193_ _06910_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14690_ VPWR VGND VPWR VGND _09671_ _09800_ _09106_ _09651_ _10157_ sky130_fd_sc_hd__a22o_2
XFILLER_0_19_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23888_ VGND VPWR VPWR VGND clk _00381_ reset_n keymem.key_mem\[13\]\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_170_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13641_ VGND VPWR _09113_ _09112_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25627_ VGND VPWR VPWR VGND clk _02120_ reset_n keymem.key_mem\[0\]\[84\] sky130_fd_sc_hd__dfrtp_2
X_22839_ VPWR VGND _06868_ keymem.rcon_logic.tmp_rcon\[0\] keymem.rcon_reg\[2\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_131_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_545 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_78_180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_168_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_196_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16360_ VGND VPWR VGND VPWR _02522_ _02520_ _02523_ _02521_ sky130_fd_sc_hd__nand3_2
X_13572_ VGND VPWR _09044_ _08982_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25558_ VGND VPWR VPWR VGND clk _02051_ reset_n keymem.key_mem\[0\]\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_195_196 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15311_ VGND VPWR VGND VPWR _10772_ _10472_ _10771_ _10751_ _10773_ sky130_fd_sc_hd__a2bb2o_2
X_12523_ VGND VPWR VGND VPWR _07786_ keymem.key_mem\[10\]\[37\] _08086_ _08088_ _08089_
+ _08069_ sky130_fd_sc_hd__a2111o_2
X_24509_ VGND VPWR VPWR VGND clk _01002_ reset_n keymem.key_mem\[9\]\[118\] sky130_fd_sc_hd__dfrtp_2
X_16291_ VPWR VGND VGND VPWR _11323_ _11280_ _11303_ _02455_ sky130_fd_sc_hd__nor3_2
XFILLER_0_26_228 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_140_1_Left_407 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25489_ VGND VPWR VPWR VGND clk _01982_ reset_n keymem.key_mem\[1\]\[74\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15242_ VPWR VGND VPWR VGND _10478_ _10541_ _10575_ _10472_ _10562_ _10705_ sky130_fd_sc_hd__a221o_2
X_18030_ VGND VPWR _03952_ _03947_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_87_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12454_ VGND VPWR enc_block.round_key\[30\] _08026_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15173_ VGND VPWR VGND VPWR _10637_ _10530_ _10604_ _10496_ _10633_ _10636_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_78_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12385_ VGND VPWR _07963_ _07632_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_111_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_151_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14124_ VPWR VGND VGND VPWR _09268_ _09293_ _09595_ _09332_ _09348_ sky130_fd_sc_hd__o22ai_2
X_19981_ VGND VPWR _00770_ _05406_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_22_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18932_ VPWR VGND VPWR VGND _04769_ _04664_ _04768_ enc_block.block_w2_reg\[18\]
+ _04709_ _00358_ sky130_fd_sc_hd__a221o_2
X_14055_ VGND VPWR VGND VPWR _09505_ keymem.prev_key1_reg\[96\] _09527_ _09429_ sky130_fd_sc_hd__nand3_2
XFILLER_0_254_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13006_ VPWR VGND VPWR VGND _08524_ keymem.key_mem\[11\]\[84\] _07809_ keymem.key_mem\[2\]\[84\]
+ _07698_ _08525_ sky130_fd_sc_hd__a221o_2
XFILLER_0_20_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_702 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18863_ VPWR VGND VGND VPWR _04654_ _04708_ _04107_ sky130_fd_sc_hd__nor2_2
XFILLER_0_24_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17814_ VGND VPWR VPWR VGND _03777_ _03804_ keymem.prev_key0_reg\[64\] _03805_ sky130_fd_sc_hd__mux2_2
XFILLER_0_197_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18794_ VGND VPWR VGND VPWR _04644_ _03951_ _04645_ _00344_ sky130_fd_sc_hd__a21o_2
XFILLER_0_238_1142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_238_1175 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17745_ VGND VPWR VPWR VGND _03719_ key[167] keymem.prev_key1_reg\[39\] _03761_ sky130_fd_sc_hd__mux2_2
X_14957_ VGND VPWR VGND VPWR _10421_ enc_block.sword_ctr_reg\[0\] enc_block.block_w1_reg\[13\]
+ enc_block.sword_ctr_reg\[1\] sky130_fd_sc_hd__and3b_2
XFILLER_0_37_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1028 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13908_ VGND VPWR _09380_ _09379_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17676_ VGND VPWR VPWR VGND _03703_ _03713_ keymem.prev_key0_reg\[17\] _03714_ sky130_fd_sc_hd__mux2_2
X_14888_ VGND VPWR VGND VPWR _09229_ _09190_ _09042_ _09666_ _10353_ sky130_fd_sc_hd__a31o_2
X_19415_ VGND VPWR VPWR VGND _05092_ _04889_ keymem.key_mem\[12\]\[7\] _05104_ sky130_fd_sc_hd__mux2_2
XFILLER_0_186_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16627_ _02780_ _02783_ _02779_ _02781_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_13839_ VGND VPWR _09311_ _09310_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_9_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_57_342 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_134_1195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_31_1112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_35_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19346_ VPWR VGND keymem.key_mem_we _05058_ _03567_ VPWR VGND sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_72_1_Left_339 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16558_ VPWR VGND VGND VPWR _09732_ _02717_ key[153] sky130_fd_sc_hd__nor2_2
XFILLER_0_174_347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15509_ VGND VPWR _10969_ keymem.prev_key1_reg\[76\] _10968_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_19277_ VPWR VGND keymem.key_mem_we _05013_ _03401_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16489_ VPWR VGND _02650_ keymem.prev_key1_reg\[55\] keymem.prev_key1_reg\[23\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_31_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18228_ VGND VPWR VPWR VGND _03973_ enc_block.block_w0_reg\[14\] _04135_ _04136_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_14_913 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_186_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_150_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_165_2_Left_636 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_667 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_108_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18159_ VGND VPWR _04073_ _08940_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21170_ VGND VPWR _01327_ _06038_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_145_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20121_ VGND VPWR _00837_ _05479_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_229_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_1230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_86 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_106_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20052_ VGND VPWR _00804_ _05443_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_42_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_830 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_225_521 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_225_532 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24860_ VGND VPWR VPWR VGND clk _01353_ reset_n keymem.key_mem\[6\]\[85\] sky130_fd_sc_hd__dfrtp_2
X_23811_ VGND VPWR VPWR VGND clk _00304_ reset_n enc_block.block_w0_reg\[30\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24791_ VGND VPWR VPWR VGND clk _01284_ reset_n keymem.key_mem\[6\]\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_197_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23742_ keymem.prev_key0_reg\[98\] clk _00239_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20954_ VGND VPWR VPWR VGND _05912_ _05010_ keymem.key_mem\[7\]\[86\] _05924_ sky130_fd_sc_hd__mux2_2
XFILLER_0_177_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_230_1415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23673_ keymem.prev_key0_reg\[29\] clk _00170_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20885_ VGND VPWR VGND VPWR _05887_ keymem.key_mem_we _03083_ _05864_ _01193_ sky130_fd_sc_hd__a31o_2
XFILLER_0_113_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25412_ VGND VPWR VPWR VGND clk _01905_ reset_n keymem.key_mem\[2\]\[125\] sky130_fd_sc_hd__dfrtp_2
X_22624_ VGND VPWR VPWR VGND _06779_ keymem.key_mem\[0\]\[2\] _09862_ _06782_ sky130_fd_sc_hd__mux2_2
XFILLER_0_152_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25343_ VGND VPWR VPWR VGND clk _01836_ reset_n keymem.key_mem\[2\]\[56\] sky130_fd_sc_hd__dfrtp_2
X_22555_ VGND VPWR VPWR VGND _06750_ keymem.key_mem\[1\]\[80\] _03330_ _06763_ sky130_fd_sc_hd__mux2_2
XFILLER_0_10_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_559 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_97_2_Left_568 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21506_ VGND VPWR VPWR VGND _06209_ _03417_ keymem.key_mem\[5\]\[90\] _06216_ sky130_fd_sc_hd__mux2_2
XFILLER_0_1_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25274_ VGND VPWR VPWR VGND clk _01767_ reset_n keymem.key_mem\[3\]\[115\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_84_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22486_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[38\] _06707_ _06706_ _04931_ _01946_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_88_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_570 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1_1098 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_133_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24225_ VGND VPWR VPWR VGND clk _00718_ reset_n keymem.key_mem\[11\]\[90\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_90_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21437_ VGND VPWR VPWR VGND _06173_ _03118_ keymem.key_mem\[5\]\[57\] _06180_ sky130_fd_sc_hd__mux2_2
XFILLER_0_43_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12170_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[8\] _07536_ _07764_ _07755_ _07765_
+ sky130_fd_sc_hd__o22a_2
X_24156_ VGND VPWR VPWR VGND clk _00649_ reset_n keymem.key_mem\[11\]\[21\] sky130_fd_sc_hd__dfrtp_2
X_21368_ VGND VPWR VPWR VGND _06140_ _02688_ keymem.key_mem\[5\]\[24\] _06144_ sky130_fd_sc_hd__mux2_2
XFILLER_0_124_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_163_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23107_ VGND VPWR VGND VPWR _03456_ _06928_ _03458_ _07031_ sky130_fd_sc_hd__a21o_2
X_20319_ VGND VPWR _00929_ _05585_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24087_ VGND VPWR VPWR VGND clk _00580_ reset_n keymem.key_mem\[12\]\[80\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_247_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21299_ VGND VPWR VPWR VGND _06098_ _03627_ keymem.key_mem\[6\]\[121\] _06106_ sky130_fd_sc_hd__mux2_2
X_23038_ VGND VPWR _02244_ _06989_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_120_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_1_Right_684 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_95_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_262_148 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15860_ VGND VPWR _11316_ _11249_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_565 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_95_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14811_ VPWR VGND VGND VPWR _10277_ _10275_ _10276_ sky130_fd_sc_hd__nand2_2
X_15791_ VGND VPWR _11247_ _11243_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_216_598 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24989_ VGND VPWR VPWR VGND clk _01482_ reset_n keymem.key_mem\[5\]\[86\] sky130_fd_sc_hd__dfrtp_2
X_17530_ VPWR VGND VGND VPWR _03597_ _02486_ _02487_ sky130_fd_sc_hd__nand2_2
X_14742_ VGND VPWR VGND VPWR _09154_ _09149_ _09204_ _09114_ _10208_ sky130_fd_sc_hd__o22a_2
XFILLER_0_98_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11954_ VGND VPWR _07557_ _07556_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_54_1123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_168_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14673_ VGND VPWR VGND VPWR _10127_ _10139_ _10140_ _10120_ _10134_ sky130_fd_sc_hd__nor4_2
X_17461_ VPWR VGND VPWR VGND _03537_ _09534_ _02979_ key[235] _03211_ _03538_ sky130_fd_sc_hd__a221o_2
XFILLER_0_135_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_170_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11885_ VGND VPWR result[109] _07506_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_104_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19200_ VGND VPWR VGND VPWR _04966_ keymem.key_mem_we _03119_ _04924_ _00429_ sky130_fd_sc_hd__a31o_2
XFILLER_0_211_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16412_ VPWR VGND VGND VPWR _11218_ _11210_ _02574_ _11205_ _11372_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_32_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13624_ VPWR VGND VPWR VGND _09031_ _09027_ _08970_ _09008_ _09096_ sky130_fd_sc_hd__or4_2
XFILLER_0_170_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17392_ VGND VPWR VGND VPWR _03478_ _09721_ _09795_ key[98] sky130_fd_sc_hd__o21a_2
XFILLER_0_131_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19131_ VPWR VGND keymem.key_mem_we _04922_ _02883_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16343_ VGND VPWR VGND VPWR _11517_ _02504_ _02506_ _02505_ sky130_fd_sc_hd__nand3_2
X_13555_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[0\] _08956_ _09027_ _08943_ _09025_
+ _09026_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_27_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12506_ VGND VPWR VGND VPWR _08074_ _07731_ keymem.key_mem\[13\]\[35\] _08071_ _08073_
+ sky130_fd_sc_hd__a211o_2
X_16274_ VPWR VGND VGND VPWR _11262_ _11305_ _02438_ _11361_ _11329_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_42_507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19062_ VGND VPWR VGND VPWR _04883_ keymem.key_mem_we _09862_ _04878_ _00374_ sky130_fd_sc_hd__a31o_2
X_13486_ VGND VPWR _08958_ _08957_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15225_ VPWR VGND VGND VPWR _10485_ _10646_ _10688_ _10521_ _10546_ sky130_fd_sc_hd__o22ai_2
X_18013_ VGND VPWR VGND VPWR _03730_ keymem.prev_key0_reg\[127\] _03940_ _03666_ _00268_
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_246_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12437_ VGND VPWR _08011_ _07761_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_22_220 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_124_299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15156_ VGND VPWR VGND VPWR _10527_ _10504_ _10545_ _10619_ _10590_ _10620_ sky130_fd_sc_hd__o32a_2
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_239_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12368_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[23\] _07577_ keymem.key_mem\[1\]\[23\]
+ _07556_ _07948_ sky130_fd_sc_hd__a22o_2
XFILLER_0_196_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14107_ VGND VPWR VGND VPWR _09578_ _09392_ _09358_ _09576_ _09333_ _09577_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_181_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15087_ VPWR VGND VPWR VGND _10550_ _10551_ _10537_ _10542_ sky130_fd_sc_hd__or3b_2
XFILLER_0_103_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19964_ VGND VPWR VPWR VGND _05389_ _10369_ keymem.key_mem\[10\]\[7\] _05397_ sky130_fd_sc_hd__mux2_2
X_12299_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[18\] _07761_ keymem.key_mem\[10\]\[18\]
+ _07674_ _07884_ sky130_fd_sc_hd__a22o_2
XFILLER_0_43_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_142_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18915_ VGND VPWR _04754_ enc_block.block_w2_reg\[25\] _04753_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_14038_ VPWR VGND VGND VPWR keymem.round_ctr_reg\[2\] keymem.round_ctr_reg\[3\] _08925_
+ _09510_ sky130_fd_sc_hd__nor3_2
XFILLER_0_103_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_638 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19895_ VGND VPWR VPWR VGND _05350_ keymem.key_mem\[11\]\[104\] _03518_ _05359_ sky130_fd_sc_hd__mux2_2
XFILLER_0_38_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_180_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18846_ VGND VPWR _04692_ enc_block.block_w0_reg\[9\] _04615_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_1172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18777_ VPWR VGND VGND VPWR _04630_ _04625_ _04628_ sky130_fd_sc_hd__nand2_2
XFILLER_0_145_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_253_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15989_ VGND VPWR VGND VPWR _11442_ _11444_ _11159_ _11158_ keylen _11445_ sky130_fd_sc_hd__o32a_2
XFILLER_0_54_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17728_ VPWR VGND VGND VPWR _03751_ _03752_ _03731_ sky130_fd_sc_hd__nor2_2
XFILLER_0_210_719 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_216_1270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_159_130 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17659_ VGND VPWR VGND VPWR _10971_ keymem.prev_key1_reg\[12\] _03702_ _03670_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_153_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_58_640 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_114_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20670_ VGND VPWR VPWR VGND _05761_ _03364_ keymem.key_mem\[8\]\[84\] _05770_ sky130_fd_sc_hd__mux2_2
XFILLER_0_70_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_110_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_312 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_50_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19329_ VGND VPWR VPWR VGND _05046_ _05045_ keymem.key_mem\[13\]\[106\] _05047_ sky130_fd_sc_hd__mux2_2
XFILLER_0_161_76 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_910 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_70_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22340_ VGND VPWR _01875_ _06660_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_264_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_954 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22271_ VGND VPWR _01842_ _06624_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_264_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_258_900 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24010_ VGND VPWR VPWR VGND clk _00503_ reset_n keymem.key_mem\[12\]\[3\] sky130_fd_sc_hd__dfrtp_2
X_21222_ VGND VPWR VPWR VGND _06065_ _03364_ keymem.key_mem\[6\]\[84\] _06066_ sky130_fd_sc_hd__mux2_2
XFILLER_0_79_83 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21153_ VGND VPWR VPWR VGND _06029_ _03067_ keymem.key_mem\[6\]\[51\] _06030_ sky130_fd_sc_hd__mux2_2
XFILLER_0_121_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20104_ VGND VPWR VPWR VGND _05469_ _03268_ keymem.key_mem\[10\]\[73\] _05471_ sky130_fd_sc_hd__mux2_2
XFILLER_0_121_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_638 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21084_ VGND VPWR _01286_ _05993_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_10_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_258_1359 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20035_ VGND VPWR _00796_ _05434_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24912_ VGND VPWR VPWR VGND clk _01405_ reset_n keymem.key_mem\[5\]\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_226_863 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24843_ VGND VPWR VPWR VGND clk _01336_ reset_n keymem.key_mem\[6\]\[68\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_213_524 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24774_ VGND VPWR VPWR VGND clk _01267_ reset_n keymem.key_mem\[7\]\[127\] sky130_fd_sc_hd__dfrtp_2
X_21986_ VPWR VGND keymem.key_mem\[3\]\[57\] _06473_ _06469_ VPWR VGND sky130_fd_sc_hd__and2_2
X_23725_ keymem.prev_key0_reg\[81\] clk _00222_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20937_ VGND VPWR VPWR VGND _05912_ _04997_ keymem.key_mem\[7\]\[78\] _05915_ sky130_fd_sc_hd__mux2_2
X_11670_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[2\] dec_new_block\[2\]
+ _07399_ sky130_fd_sc_hd__mux2_2
X_23656_ keymem.prev_key0_reg\[12\] clk _00153_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20868_ VGND VPWR VPWR VGND _05867_ _04947_ keymem.key_mem\[7\]\[46\] _05878_ sky130_fd_sc_hd__mux2_2
X_22607_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[117\] _06777_ _06776_ _05069_ _02025_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_14_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23587_ VGND VPWR VPWR VGND clk _00088_ reset_n keymem.key_mem\[14\]\[76\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_265_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20799_ VPWR VGND keymem.key_mem\[7\]\[14\] _05841_ _05830_ VPWR VGND sky130_fd_sc_hd__and2_2
X_25326_ VGND VPWR VPWR VGND clk _01819_ reset_n keymem.key_mem\[2\]\[39\] sky130_fd_sc_hd__dfrtp_2
X_13340_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[117\] _07924_ keymem.key_mem\[8\]\[117\]
+ _07878_ _08826_ sky130_fd_sc_hd__a22o_2
XFILLER_0_146_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22538_ VGND VPWR _06757_ _03227_ _01976_ _06756_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_8_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25257_ VGND VPWR VPWR VGND clk _01750_ reset_n keymem.key_mem\[3\]\[98\] sky130_fd_sc_hd__dfrtp_2
X_13271_ VGND VPWR VGND VPWR _07839_ keymem.key_mem\[11\]\[110\] _08761_ _08763_ _08764_
+ _07574_ sky130_fd_sc_hd__a2111o_2
X_22469_ VGND VPWR VPWR VGND _06726_ keymem.key_mem\[1\]\[28\] _02787_ _06729_ sky130_fd_sc_hd__mux2_2
XFILLER_0_161_361 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_106_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15010_ VPWR VGND VGND VPWR _10473_ _10474_ _10472_ sky130_fd_sc_hd__nor2_2
XFILLER_0_121_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24208_ VGND VPWR VPWR VGND clk _00701_ reset_n keymem.key_mem\[11\]\[73\] sky130_fd_sc_hd__dfrtp_2
X_12222_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[12\] _07812_ keymem.key_mem\[1\]\[12\]
+ _07714_ _07813_ sky130_fd_sc_hd__a22o_2
XFILLER_0_66_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25188_ VGND VPWR VPWR VGND clk _01681_ reset_n keymem.key_mem\[3\]\[29\] sky130_fd_sc_hd__dfrtp_2
X_12153_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[7\] _07748_ keymem.key_mem\[12\]\[7\]
+ _07722_ _07749_ sky130_fd_sc_hd__a22o_2
X_24139_ VGND VPWR VPWR VGND clk _00632_ reset_n keymem.key_mem\[11\]\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16961_ VGND VPWR _03091_ _03090_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12084_ VGND VPWR _07683_ _07595_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18700_ VGND VPWR _04560_ _03981_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15912_ VPWR VGND VGND VPWR _11367_ _11368_ _11303_ sky130_fd_sc_hd__nor2_2
XFILLER_0_159_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19680_ VGND VPWR _05246_ _05242_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16892_ VGND VPWR VPWR VGND _11160_ _11441_ _02864_ _03028_ sky130_fd_sc_hd__or3_2
XFILLER_0_95_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_84_1_Right_685 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_246_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18631_ VGND VPWR _04499_ _04497_ _04498_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_159_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15843_ VPWR VGND VGND VPWR _11293_ _11296_ _11298_ _11292_ _11299_ sky130_fd_sc_hd__and4b_2
XFILLER_0_95_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18562_ VPWR VGND VGND VPWR _04437_ _04434_ _04436_ sky130_fd_sc_hd__nand2_2
X_15774_ VGND VPWR VGND VPWR _11230_ _11229_ _11228_ _11227_ _11226_ sky130_fd_sc_hd__and4_2
X_12986_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[82\] _08125_ keymem.key_mem\[8\]\[82\]
+ _07958_ _08507_ sky130_fd_sc_hd__a22o_2
XFILLER_0_188_247 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_59_415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_231_1009 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17513_ VGND VPWR VGND VPWR _03582_ _10328_ _02877_ key[115] sky130_fd_sc_hd__o21a_2
XFILLER_0_8_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14725_ VGND VPWR VPWR VGND _09796_ key[5] _10192_ _10191_ _10188_ sky130_fd_sc_hd__o211a_2
X_18493_ VPWR VGND VGND VPWR _04375_ _04372_ _04374_ sky130_fd_sc_hd__nand2_2
XFILLER_0_262_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11937_ VGND VPWR _07540_ _07539_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_200_752 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17444_ VGND VPWR VPWR VGND _10378_ _03522_ key[233] _03523_ sky130_fd_sc_hd__mux2_2
X_14656_ VGND VPWR VPWR VGND _10121_ _10122_ _09591_ _10123_ sky130_fd_sc_hd__or3_2
X_11868_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[5\] dec_new_block\[101\]
+ _07498_ sky130_fd_sc_hd__mux2_2
XFILLER_0_262_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13607_ VPWR VGND VPWR VGND _09014_ _09015_ _09045_ _09043_ _09079_ sky130_fd_sc_hd__or4_2
XFILLER_0_7_729 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17375_ VGND VPWR VGND VPWR _09527_ _09526_ _03463_ _10092_ sky130_fd_sc_hd__a21oi_2
X_11799_ VGND VPWR result[66] _07463_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14587_ VPWR VGND VPWR VGND _10053_ _10054_ _10055_ _10048_ _10051_ sky130_fd_sc_hd__or4b_2
XFILLER_0_32_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19114_ VGND VPWR VGND VPWR _04912_ keymem.key_mem_we _02721_ _04908_ _00397_ sky130_fd_sc_hd__a31o_2
XFILLER_0_171_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_54_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16326_ VGND VPWR VGND VPWR _02487_ _02486_ _02489_ _02484_ sky130_fd_sc_hd__a21oi_2
X_13538_ VGND VPWR _09010_ _08963_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_171_136 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_166_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19045_ VGND VPWR _04870_ _04667_ _04869_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16257_ VGND VPWR VGND VPWR _02419_ _02418_ _11563_ _02347_ _02421_ _02420_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_28_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13469_ VPWR VGND VGND VPWR _08940_ _08941_ _08938_ sky130_fd_sc_hd__nor2_2
XFILLER_0_2_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15208_ VPWR VGND VGND VPWR _10671_ _10669_ _10670_ sky130_fd_sc_hd__nand2_2
X_16188_ VGND VPWR VGND VPWR _11210_ _11241_ _11482_ _11275_ _02353_ sky130_fd_sc_hd__o22a_2
XFILLER_0_2_489 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_11_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15139_ VPWR VGND VPWR VGND _10457_ _10435_ _10444_ _10443_ _10603_ sky130_fd_sc_hd__or4_2
XFILLER_0_11_779 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_103_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19947_ VGND VPWR _05387_ _05386_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_103_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_10 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19878_ VGND VPWR _05350_ _05242_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_78_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_138_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_177_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18829_ VPWR VGND VPWR VGND _04677_ _04603_ _04675_ sky130_fd_sc_hd__or2_2
XFILLER_0_74_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_39_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21840_ VGND VPWR _01643_ _06392_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_223_888 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_222_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_250_696 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_253_1289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_210_527 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21771_ VGND VPWR _01610_ _06356_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23510_ VGND VPWR VPWR VGND clk _00006_ reset_n aes_core_ctrl_reg\[2\] sky130_fd_sc_hd__dfrtp_2
X_20722_ VGND VPWR _01120_ _05797_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24490_ VGND VPWR VPWR VGND clk _00983_ reset_n keymem.key_mem\[9\]\[99\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_114_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_2_Left_580 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_188_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23441_ VPWR VGND VPWR VGND _07307_ _04065_ enc_block.block_w3_reg\[24\] _03953_
+ _07308_ sky130_fd_sc_hd__a22o_2
XFILLER_0_110_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20653_ VGND VPWR _05761_ _05679_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_11_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23372_ VGND VPWR _07246_ enc_block.block_w0_reg\[16\] enc_block.block_w0_reg\[23\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20584_ VGND VPWR _05725_ _05679_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_184_1339 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_149_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_315 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_264_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25111_ VGND VPWR VPWR VGND clk _01604_ reset_n keymem.key_mem\[4\]\[80\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_150_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_646 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_85_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22323_ VGND VPWR _01867_ _06651_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_46_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_860 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_103_214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_264_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25042_ VGND VPWR VPWR VGND clk _01535_ reset_n keymem.key_mem\[4\]\[11\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22254_ VGND VPWR _01834_ _06615_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_42_882 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_108_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_595 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21205_ VGND VPWR VPWR VGND _06052_ _03295_ keymem.key_mem\[6\]\[76\] _06057_ sky130_fd_sc_hd__mux2_2
X_22185_ VGND VPWR _01801_ _06579_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_121_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21136_ VGND VPWR VPWR VGND _06018_ _02985_ keymem.key_mem\[6\]\[43\] _06021_ sky130_fd_sc_hd__mux2_2
XFILLER_0_121_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21067_ VGND VPWR _01278_ _05984_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_201_1391 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20018_ VGND VPWR VPWR VGND _05424_ _02873_ keymem.key_mem\[10\]\[32\] _05426_ sky130_fd_sc_hd__mux2_2
XFILLER_0_195_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_226_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_216_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_57_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12840_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[67\] _07644_ _08375_ _08371_ _08376_
+ sky130_fd_sc_hd__o22a_2
X_24826_ VGND VPWR VPWR VGND clk _01319_ reset_n keymem.key_mem\[6\]\[51\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_236_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_201_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12771_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[60\] _08259_ _08313_ _08309_ _08314_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_240_173 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_198_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21969_ VGND VPWR VPWR VGND _06462_ _04953_ keymem.key_mem\[3\]\[49\] _06464_ sky130_fd_sc_hd__mux2_2
X_24757_ VGND VPWR VPWR VGND clk _01250_ reset_n keymem.key_mem\[7\]\[110\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_51_1115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11722_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[28\] dec_new_block\[28\]
+ _07425_ sky130_fd_sc_hd__mux2_2
X_14510_ VPWR VGND VGND VPWR _09141_ _09097_ _09114_ _09658_ _09979_ _09978_ sky130_fd_sc_hd__o221a_2
X_15490_ VGND VPWR _10949_ _10553_ _10950_ _10856_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_28_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23708_ keymem.prev_key0_reg\[64\] clk _00205_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_56_429 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24688_ VGND VPWR VPWR VGND clk _01181_ reset_n keymem.key_mem\[7\]\[41\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_132_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14441_ VPWR VGND VGND VPWR _09411_ _09910_ _09426_ sky130_fd_sc_hd__nor2_2
X_11653_ VGND VPWR VGND VPWR _00010_ keymem.key_mem_we _07384_ _07383_ _07389_ keymem.round_ctr_rst
+ sky130_fd_sc_hd__a41o_2
X_23639_ VPWR VGND VPWR VGND ready reset_n _00140_ clk sky130_fd_sc_hd__dfstp_2
XFILLER_0_232_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_167_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_153_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14372_ _09086_ _09842_ _09047_ _09199_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_17160_ _10817_ _03270_ keymem.prev_key0_reg\[74\] _10818_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_64_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_175 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_167_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16111_ _11396_ _11565_ _11224_ _11292_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_247_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13323_ VGND VPWR VGND VPWR _08811_ _07839_ keymem.key_mem\[11\]\[115\] _08808_ _08810_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_153_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25309_ VGND VPWR VPWR VGND clk _01802_ reset_n keymem.key_mem\[2\]\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_64_1509 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17091_ VPWR VGND VPWR VGND _03208_ _02497_ _03204_ key[194] _03027_ _03209_ sky130_fd_sc_hd__a221o_2
XFILLER_0_51_145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16042_ VGND VPWR VGND VPWR _11497_ _11221_ _11286_ _11167_ _11174_ sky130_fd_sc_hd__a211o_2
X_13254_ VPWR VGND VPWR VGND _08748_ keymem.key_mem\[13\]\[108\] _08125_ keymem.key_mem\[4\]\[108\]
+ _07854_ _08749_ sky130_fd_sc_hd__a221o_2
XFILLER_0_33_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_243_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12205_ VPWR VGND VPWR VGND _07796_ keymem.key_mem\[10\]\[11\] _07742_ keymem.key_mem\[4\]\[11\]
+ _07692_ _07797_ sky130_fd_sc_hd__a221o_2
XFILLER_0_86_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13185_ VGND VPWR enc_block.round_key\[101\] _08686_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_161_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19801_ VGND VPWR VPWR VGND _05303_ keymem.key_mem\[11\]\[59\] _03140_ _05310_ sky130_fd_sc_hd__mux2_2
XFILLER_0_249_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_104_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12136_ VGND VPWR _07732_ _07545_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17993_ VGND VPWR VGND VPWR _02647_ keymem.prev_key1_reg\[121\] _03679_ _03927_ sky130_fd_sc_hd__a21o_2
XFILLER_0_100_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19732_ VGND VPWR VPWR VGND _05270_ keymem.key_mem\[11\]\[26\] _02743_ _05274_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_81_1_Left_348 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_252_917 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16944_ VGND VPWR VPWR VGND _02986_ keymem.key_mem\[14\]\[52\] _03075_ _03076_ sky130_fd_sc_hd__mux2_2
XFILLER_0_236_468 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12067_ VGND VPWR _07667_ _07586_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_223_118 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_174_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19663_ VGND VPWR _00623_ _05235_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16875_ VPWR VGND VGND VPWR keylen _03012_ keymem.prev_key1_reg\[46\] _10287_ _11048_
+ _03013_ sky130_fd_sc_hd__a311o_2
XFILLER_0_126_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_254_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_1_Right_686 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18614_ VPWR VGND VPWR VGND _04483_ block[82] _04330_ enc_block.block_w2_reg\[18\]
+ _04425_ _04484_ sky130_fd_sc_hd__a221o_2
XFILLER_0_215_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_204_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15826_ VGND VPWR _11282_ _11281_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_56_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19594_ VGND VPWR VGND VPWR _05199_ keymem.key_mem_we _03418_ _05187_ _00590_ sky130_fd_sc_hd__a31o_2
XPHY_EDGE_ROW_174_2_Left_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_250_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18545_ VPWR VGND _04422_ _04421_ enc_block.round_key\[75\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15757_ VGND VPWR VGND VPWR _11213_ enc_block.block_w2_reg\[16\] enc_block.sword_ctr_reg\[1\]
+ enc_block.sword_ctr_reg\[0\] sky130_fd_sc_hd__and3b_2
XFILLER_0_59_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12969_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[80\] _07577_ keymem.key_mem\[4\]\[80\]
+ _07550_ _08492_ sky130_fd_sc_hd__a22o_2
XFILLER_0_143_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14708_ VGND VPWR VGND VPWR _09234_ _10173_ _10174_ _09944_ _09106_ _10175_ sky130_fd_sc_hd__o41a_2
X_18476_ VPWR VGND VPWR VGND _04359_ block[68] _04351_ enc_block.block_w0_reg\[4\]
+ _03954_ _04360_ sky130_fd_sc_hd__a221o_2
XFILLER_0_111_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15688_ VGND VPWR VGND VPWR _11144_ _11109_ _11145_ _11111_ sky130_fd_sc_hd__nand3_2
XFILLER_0_150_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17427_ VPWR VGND VGND VPWR _03508_ key[231] _03077_ sky130_fd_sc_hd__nand2_2
X_14639_ VPWR VGND VGND VPWR _09487_ _09350_ _09423_ _09456_ _10106_ _10105_ sky130_fd_sc_hd__o221a_2
XFILLER_0_74_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_111_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_74_259 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_43_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_462 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17358_ VGND VPWR VGND VPWR _11624_ _03446_ _02817_ _02822_ _03448_ sky130_fd_sc_hd__a31o_2
XFILLER_0_132_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16309_ VGND VPWR VGND VPWR _02471_ _02470_ _02473_ _02472_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_125_350 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17289_ VGND VPWR VGND VPWR _02708_ key[215] _03386_ _02656_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_261_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19028_ VGND VPWR _04855_ enc_block.block_w3_reg\[20\] _04854_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_222_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23990_ VGND VPWR VPWR VGND clk _00483_ reset_n keymem.key_mem\[13\]\[111\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_255_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_991 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22941_ VGND VPWR _02204_ _06932_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_78_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1224 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_223_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_207_192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22872_ VGND VPWR _06888_ _06878_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25660_ VGND VPWR VPWR VGND clk _02153_ reset_n keymem.key_mem\[0\]\[117\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24611_ VGND VPWR VPWR VGND clk _01104_ reset_n keymem.key_mem\[8\]\[92\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_218_1195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21823_ VGND VPWR _01635_ _06383_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_6_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25591_ VGND VPWR VPWR VGND clk _02084_ reset_n keymem.key_mem\[0\]\[48\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_214_1037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_210_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1376 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_211_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24542_ VGND VPWR VPWR VGND clk _01035_ reset_n keymem.key_mem\[8\]\[23\] sky130_fd_sc_hd__dfrtp_2
X_21754_ VGND VPWR _01602_ _06347_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_114_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20705_ VGND VPWR _01112_ _05788_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24473_ VGND VPWR VPWR VGND clk _00966_ reset_n keymem.key_mem\[9\]\[82\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_175_261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21685_ VGND VPWR _01569_ _06311_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_11_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23424_ VPWR VGND VPWR VGND _07292_ _04064_ enc_block.block_w0_reg\[22\] _03952_
+ _07293_ sky130_fd_sc_hd__a22o_2
XFILLER_0_149_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20636_ VGND VPWR _01079_ _05752_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_85_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_18_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23355_ VPWR VGND _07231_ enc_block.block_w1_reg\[14\] enc_block.block_w2_reg\[6\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_61_443 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20567_ VGND VPWR _01046_ _05716_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_85_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1217 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22306_ VGND VPWR _01859_ _06642_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_131_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23286_ VPWR VGND VPWR VGND _07169_ _07166_ _07168_ sky130_fd_sc_hd__or2_2
XFILLER_0_143_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20498_ VGND VPWR _05680_ _05679_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25025_ VGND VPWR VPWR VGND clk _01518_ reset_n keymem.key_mem\[5\]\[122\] sky130_fd_sc_hd__dfrtp_2
X_22237_ VGND VPWR _01826_ _06606_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_246_711 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_896 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22168_ VGND VPWR _01793_ _06570_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21119_ VGND VPWR VPWR VGND _06007_ _02903_ keymem.key_mem\[6\]\[35\] _06012_ sky130_fd_sc_hd__mux2_2
XFILLER_0_246_777 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14990_ VGND VPWR VPWR VGND _10453_ _10409_ _10451_ _10454_ sky130_fd_sc_hd__or3_2
XFILLER_0_22_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22099_ VGND VPWR _01762_ _06532_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_261_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13941_ VGND VPWR VGND VPWR _09302_ _09397_ _09336_ _09404_ _09413_ sky130_fd_sc_hd__o22a_2
XFILLER_0_96_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16660_ VGND VPWR VGND VPWR keymem.rcon_logic.tmp_rcon\[7\] _02572_ _02814_ _02586_
+ sky130_fd_sc_hd__a21bo_2
X_13872_ VGND VPWR VGND VPWR _09333_ _09336_ _09343_ _09341_ _09344_ sky130_fd_sc_hd__o22a_2
XFILLER_0_57_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_353 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15611_ VPWR VGND VGND VPWR _10593_ _10639_ _10535_ _10543_ _11069_ _10555_ sky130_fd_sc_hd__o221a_2
X_12823_ VGND VPWR VGND VPWR _08360_ _07841_ keymem.key_mem\[4\]\[66\] _08359_ _07896_
+ sky130_fd_sc_hd__a211o_2
X_24809_ VGND VPWR VPWR VGND clk _01302_ reset_n keymem.key_mem\[6\]\[34\] sky130_fd_sc_hd__dfrtp_2
X_16591_ VGND VPWR VGND VPWR _09923_ _09883_ _02748_ _09240_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_201_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25789_ keymem.prev_key1_reg\[105\] clk _02282_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_158_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18330_ VPWR VGND VGND VPWR _04228_ _04229_ _04077_ sky130_fd_sc_hd__nor2_2
X_15542_ VPWR VGND VPWR VGND _10778_ _11000_ _10808_ _10781_ _11001_ sky130_fd_sc_hd__or4_2
XFILLER_0_55_1092 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_738 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12754_ VPWR VGND VPWR VGND _08297_ keymem.key_mem\[9\]\[59\] _07593_ keymem.key_mem\[8\]\[59\]
+ _07753_ _08298_ sky130_fd_sc_hd__a221o_2
XFILLER_0_173_209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11705_ VGND VPWR result[19] _07416_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18261_ VGND VPWR VGND VPWR _04165_ _04164_ _04166_ _03966_ sky130_fd_sc_hd__a21oi_2
X_15473_ VPWR VGND VGND VPWR _10511_ _10933_ _10609_ sky130_fd_sc_hd__nor2_2
X_12685_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[52\] _07568_ keymem.key_mem\[2\]\[52\]
+ _07732_ _08236_ sky130_fd_sc_hd__a22o_2
XFILLER_0_56_259 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_126_114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_181_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17212_ VGND VPWR VGND VPWR _03316_ _11107_ _03317_ keylen sky130_fd_sc_hd__a21oi_2
X_14424_ VGND VPWR VGND VPWR _09893_ _09564_ _09312_ _09475_ _09392_ _09892_ sky130_fd_sc_hd__o221ai_2
X_11636_ VPWR VGND VPWR VGND _00000_ _07375_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18192_ VGND VPWR _04103_ _03955_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_4_507 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17143_ VGND VPWR VPWR VGND _02864_ _10655_ keymem.prev_key0_reg\[72\] _03255_ sky130_fd_sc_hd__or3_2
XFILLER_0_141_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14355_ VGND VPWR VGND VPWR _09095_ _09141_ _09114_ _09069_ _09825_ sky130_fd_sc_hd__o22a_2
XFILLER_0_243_1200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_68_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13306_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[114\] _07788_ keymem.key_mem\[2\]\[114\]
+ _08116_ _08795_ sky130_fd_sc_hd__a22o_2
X_14286_ VGND VPWR VPWR VGND _09468_ _09363_ _09373_ _09756_ sky130_fd_sc_hd__or3_2
XFILLER_0_243_1244 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17074_ VGND VPWR _03194_ _03193_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_97_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1217 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16025_ VGND VPWR VGND VPWR _11325_ _11298_ _11480_ _11464_ sky130_fd_sc_hd__a21oi_2
X_13237_ VPWR VGND VPWR VGND keymem.key_mem\[4\]\[107\] _07693_ keymem.key_mem\[1\]\[107\]
+ _07715_ _08733_ sky130_fd_sc_hd__a22o_2
XFILLER_0_20_340 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_582 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13168_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[100\] _07618_ keymem.key_mem\[4\]\[100\]
+ _07551_ _08671_ sky130_fd_sc_hd__a22o_2
XFILLER_0_104_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_541 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12119_ VGND VPWR _07716_ _07590_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17976_ VGND VPWR VPWR VGND _03896_ _03915_ keymem.prev_key0_reg\[115\] _03916_ sky130_fd_sc_hd__mux2_2
X_13099_ VGND VPWR VGND VPWR _07648_ keymem.key_mem\[2\]\[93\] _08606_ _08608_ _08609_
+ _08599_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_104_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19715_ VGND VPWR VPWR VGND _05259_ keymem.key_mem\[11\]\[18\] _02340_ _05265_ sky130_fd_sc_hd__mux2_2
X_16927_ VPWR VGND VPWR VGND _03060_ key[51] _08935_ sky130_fd_sc_hd__or2_2
XFILLER_0_174_1316 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_79_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_89 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_75_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19646_ VGND VPWR _00615_ _05226_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_189_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16858_ VGND VPWR VGND VPWR _02998_ _02996_ _02991_ _02990_ _02997_ sky130_fd_sc_hd__o211ai_2
XPHY_EDGE_ROW_86_1_Right_687 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_219_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15809_ VGND VPWR _11265_ _11264_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_75_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19577_ VPWR VGND keymem.key_mem\[12\]\[82\] _05191_ _05173_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_137_1182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16789_ VGND VPWR VPWR VGND _02884_ keymem.key_mem\[14\]\[38\] _02934_ _02935_ sky130_fd_sc_hd__mux2_2
X_18528_ VPWR VGND VGND VPWR _04380_ _04407_ _04086_ sky130_fd_sc_hd__nor2_2
XFILLER_0_62_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1132 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_47_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_157_250 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_30_1018 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18459_ VGND VPWR _04344_ enc_block.block_w0_reg\[7\] _04343_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_771 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21470_ VGND VPWR _01468_ _06197_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_185_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_635 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_117_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_172_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_55_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20421_ VGND VPWR VPWR VGND _05638_ _03452_ keymem.key_mem\[9\]\[94\] _05639_ sky130_fd_sc_hd__mux2_2
XFILLER_0_86_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_47_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23140_ VGND VPWR VGND VPWR _03211_ key[235] _02979_ _07052_ sky130_fd_sc_hd__a21o_2
X_20352_ VGND VPWR VPWR VGND _05602_ _03162_ keymem.key_mem\[9\]\[61\] _05603_ sky130_fd_sc_hd__mux2_2
XFILLER_0_261_1333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_226_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_830 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_113_364 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_226_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23071_ VGND VPWR _02257_ _07009_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_140_161 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20283_ VGND VPWR _00912_ _05566_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_105_1148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22022_ VGND VPWR VPWR VGND _06462_ _04989_ keymem.key_mem\[3\]\[74\] _06492_ sky130_fd_sc_hd__mux2_2
XFILLER_0_122_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_220_1052 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_196_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_243_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_157_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23973_ VGND VPWR VPWR VGND clk _00466_ reset_n keymem.key_mem\[13\]\[94\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_157_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25712_ keymem.prev_key1_reg\[28\] clk _02205_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_93_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22924_ VGND VPWR _02199_ _06920_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_233_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_460 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_39_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25643_ VGND VPWR VPWR VGND clk _02136_ reset_n keymem.key_mem\[0\]\[100\] sky130_fd_sc_hd__dfrtp_2
X_22855_ VPWR VGND VGND VPWR _06876_ keymem.round_ctr_reg\[3\] _05818_ sky130_fd_sc_hd__nand2_2
XFILLER_0_233_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21806_ VGND VPWR _01627_ _06374_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22786_ VGND VPWR VPWR VGND _06784_ keymem.key_mem\[0\]\[92\] _03435_ _06854_ sky130_fd_sc_hd__mux2_2
X_25574_ VGND VPWR VPWR VGND clk _02067_ reset_n keymem.key_mem\[0\]\[31\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_151_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21737_ VGND VPWR _01594_ _06338_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24525_ VGND VPWR VPWR VGND clk _01018_ reset_n keymem.key_mem\[8\]\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_376 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_30_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12470_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[32\] _08016_ keymem.key_mem\[6\]\[32\]
+ _07908_ _08041_ sky130_fd_sc_hd__a22o_2
XFILLER_0_4_1085 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24456_ VGND VPWR VPWR VGND clk _00949_ reset_n keymem.key_mem\[9\]\[65\] sky130_fd_sc_hd__dfrtp_2
X_21668_ VGND VPWR _01561_ _06302_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_34_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_62_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23407_ VGND VPWR _07278_ _07275_ _07277_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_123_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20619_ VGND VPWR _01071_ _05743_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24387_ VGND VPWR VPWR VGND clk _00880_ reset_n keymem.key_mem\[10\]\[124\] sky130_fd_sc_hd__dfrtp_2
X_21599_ VGND VPWR _01528_ _06266_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_62_774 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14140_ VGND VPWR VGND VPWR _09431_ _09399_ _09443_ _09363_ _09373_ _09611_ sky130_fd_sc_hd__o32a_2
XFILLER_0_61_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23338_ VGND VPWR VGND VPWR _07214_ _07213_ _07216_ _07212_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_244_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14071_ VGND VPWR _00012_ _09542_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23269_ VPWR VGND VPWR VGND _07153_ block[6] _04837_ enc_block.block_w2_reg\[6\]
+ _04798_ _07154_ sky130_fd_sc_hd__a221o_2
XFILLER_0_131_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_162_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13022_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[85\] _07645_ _08539_ _08535_ _08540_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_259_891 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25008_ VGND VPWR VPWR VGND clk _01501_ reset_n keymem.key_mem\[5\]\[105\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_197_1338 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17830_ VGND VPWR VPWR VGND _03812_ key[197] keymem.prev_key1_reg\[69\] _03816_ sky130_fd_sc_hd__mux2_2
XFILLER_0_207_906 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_101_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_238_77 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_238_1313 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_246_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17761_ VGND VPWR _00185_ _03771_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14973_ VGND VPWR _10437_ _10436_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_107_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19500_ VGND VPWR _00546_ _05149_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16712_ VGND VPWR _02864_ _09516_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13924_ VGND VPWR _09396_ _09395_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17692_ VGND VPWR _00163_ _03724_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_18_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_599 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_202_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_254_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19431_ VGND VPWR VGND VPWR _05112_ keymem.key_mem_we _11099_ _05109_ _00514_ sky130_fd_sc_hd__a31o_2
X_16643_ VGND VPWR VPWR VGND _02796_ _02691_ _02798_ _09514_ _02797_ sky130_fd_sc_hd__o211a_2
X_13855_ VGND VPWR _09327_ _09326_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_18_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12806_ VGND VPWR VGND VPWR _07737_ keymem.key_mem\[1\]\[64\] _08342_ _08344_ _08345_
+ _07574_ sky130_fd_sc_hd__a2111o_2
X_19362_ VPWR VGND keymem.key_mem_we _05069_ _03600_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_186_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16574_ VGND VPWR VPWR VGND _11109_ _02731_ key[26] _02732_ sky130_fd_sc_hd__mux2_2
X_13786_ VGND VPWR VGND VPWR enc_block.block_w1_reg\[26\] _08985_ _09022_ _09256_
+ _09258_ _09257_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_201_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_130_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18313_ VGND VPWR _04213_ _03979_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_96_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15525_ VPWR VGND VGND VPWR _10518_ _10604_ _10984_ _10510_ _10611_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_57_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_139_261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19293_ VGND VPWR _00466_ _05022_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12737_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[57\] _07594_ keymem.key_mem\[4\]\[57\]
+ _07550_ _08283_ sky130_fd_sc_hd__a22o_2
XFILLER_0_70_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_210_1243 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_719 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_84_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18244_ VGND VPWR VGND VPWR _04147_ _04150_ _03974_ _04151_ enc_block.block_w0_reg\[15\]
+ sky130_fd_sc_hd__o2bb2a_2
X_15456_ VGND VPWR _10916_ keymem.prev_key0_reg\[12\] _10915_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_12668_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[50\] _08145_ _08220_ _08215_ _08221_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_5_816 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_154_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14407_ VPWR VGND VGND VPWR _09386_ _09876_ _09330_ sky130_fd_sc_hd__nor2_2
X_18175_ VPWR VGND VPWR VGND _04087_ _04040_ _04084_ enc_block.block_w0_reg\[9\] _03976_
+ _00283_ sky130_fd_sc_hd__a221o_2
X_15387_ VGND VPWR VGND VPWR _10449_ _10476_ _10587_ _10530_ _10848_ sky130_fd_sc_hd__o22a_2
XFILLER_0_29_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_240 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12599_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[44\] _07685_ keymem.key_mem\[8\]\[44\]
+ _07654_ _08158_ sky130_fd_sc_hd__a22o_2
X_17126_ VGND VPWR _03240_ _10366_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_13_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14338_ VPWR VGND VPWR VGND _09805_ _09807_ _09808_ _09799_ _09802_ sky130_fd_sc_hd__or4b_2
XFILLER_0_68_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_424 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17057_ VPWR VGND VPWR VGND _03178_ keymem.prev_key1_reg\[63\] sky130_fd_sc_hd__inv_2
X_14269_ VPWR VGND VPWR VGND _09736_ _09738_ _09739_ _09587_ _09735_ sky130_fd_sc_hd__or4b_2
XFILLER_0_29_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16008_ VPWR VGND VGND VPWR _11463_ _11461_ _11462_ sky130_fd_sc_hd__nand2_2
XFILLER_0_141_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_110_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_139_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17959_ VGND VPWR VPWR VGND _03876_ key[238] keymem.prev_key1_reg\[110\] _03904_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_252_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20970_ VGND VPWR VPWR VGND _05912_ _05021_ keymem.key_mem\[7\]\[94\] _05932_ sky130_fd_sc_hd__mux2_2
XFILLER_0_36_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_215_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19629_ VGND VPWR VPWR VGND _05216_ _05048_ keymem.key_mem\[12\]\[107\] _05218_ sky130_fd_sc_hd__mux2_2
XFILLER_0_177_312 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_87_1_Right_688 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22640_ VGND VPWR _02044_ _06791_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_48_524 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_169_1_Left_436 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_152_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_610 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22571_ VGND VPWR VPWR VGND _06701_ keymem.key_mem\[1\]\[90\] _03418_ _06769_ sky130_fd_sc_hd__mux2_2
XFILLER_0_180_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_2_Left_608 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24310_ VGND VPWR VPWR VGND clk _00803_ reset_n keymem.key_mem\[10\]\[47\] sky130_fd_sc_hd__dfrtp_2
X_21522_ VGND VPWR _01493_ _06224_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_192_359 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25290_ VGND VPWR VPWR VGND clk _01783_ reset_n keymem.key_mem\[2\]\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_180_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_267_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_8_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24241_ VGND VPWR VPWR VGND clk _00734_ reset_n keymem.key_mem\[11\]\[106\] sky130_fd_sc_hd__dfrtp_2
X_21453_ VGND VPWR _01460_ _06188_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20404_ VGND VPWR VPWR VGND _05627_ _03383_ keymem.key_mem\[9\]\[86\] _05630_ sky130_fd_sc_hd__mux2_2
X_24172_ VGND VPWR VPWR VGND clk _00665_ reset_n keymem.key_mem\[11\]\[37\] sky130_fd_sc_hd__dfrtp_2
X_21384_ VGND VPWR _01427_ _06152_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23123_ VGND VPWR _03498_ _02919_ _07041_ _03495_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_4_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20335_ VGND VPWR VPWR VGND _05591_ _03083_ keymem.key_mem\[9\]\[53\] _05594_ sky130_fd_sc_hd__mux2_2
X_23054_ VGND VPWR _02250_ _06999_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_222_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20266_ VGND VPWR _00904_ _05557_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22005_ VGND VPWR VPWR VGND _06462_ _04977_ keymem.key_mem\[3\]\[66\] _06483_ sky130_fd_sc_hd__mux2_2
XFILLER_0_256_883 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_228_574 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20197_ VGND VPWR _00873_ _05519_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_228_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_228_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11970_ VGND VPWR _07573_ _07572_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23956_ VGND VPWR VPWR VGND clk _00449_ reset_n keymem.key_mem\[13\]\[77\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_118_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22907_ VGND VPWR VPWR VGND _06878_ _06909_ keymem.prev_key1_reg\[16\] _06910_ sky130_fd_sc_hd__mux2_2
XFILLER_0_211_430 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23887_ VGND VPWR VPWR VGND clk _00380_ reset_n keymem.key_mem\[13\]\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_975 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13640_ VPWR VGND VPWR VGND _08963_ _09027_ _09017_ _09009_ _09112_ sky130_fd_sc_hd__or4_2
X_25626_ VGND VPWR VPWR VGND clk _02119_ reset_n keymem.key_mem\[0\]\[83\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_170_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22838_ VGND VPWR VGND VPWR keymem.rcon_reg\[2\] _06862_ keymem.rcon_logic.tmp_rcon\[2\]
+ _06863_ _02166_ sky130_fd_sc_hd__o22a_2
XFILLER_0_128_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13571_ VGND VPWR _09043_ _08977_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25557_ VGND VPWR VPWR VGND clk _02050_ reset_n keymem.key_mem\[0\]\[14\] sky130_fd_sc_hd__dfrtp_2
X_22769_ VGND VPWR VPWR VGND _06833_ keymem.key_mem\[0\]\[82\] _03347_ _06847_ sky130_fd_sc_hd__mux2_2
XFILLER_0_66_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15310_ VPWR VGND VGND VPWR _10469_ _10584_ _10772_ _10563_ _10504_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_66_376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1057 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12522_ VPWR VGND VPWR VGND _08087_ keymem.key_mem\[3\]\[37\] _07844_ keymem.key_mem\[14\]\[37\]
+ _08032_ _08088_ sky130_fd_sc_hd__a221o_2
X_24508_ VGND VPWR VPWR VGND clk _01001_ reset_n keymem.key_mem\[9\]\[117\] sky130_fd_sc_hd__dfrtp_2
X_16290_ VPWR VGND VPWR VGND _02452_ _02453_ _02454_ _02450_ _02451_ sky130_fd_sc_hd__or4b_2
XFILLER_0_136_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25488_ VGND VPWR VPWR VGND clk _01981_ reset_n keymem.key_mem\[1\]\[73\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_168_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15241_ VPWR VGND VPWR VGND _10703_ _10704_ _10701_ _10702_ sky130_fd_sc_hd__or3b_2
XPHY_EDGE_ROW_90_1_Left_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24439_ VGND VPWR VPWR VGND clk _00932_ reset_n keymem.key_mem\[9\]\[48\] sky130_fd_sc_hd__dfrtp_2
X_12453_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[30\] _07793_ _08025_ _08021_ _08026_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_87_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_65_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15172_ VGND VPWR VGND VPWR _10484_ _10594_ _10540_ _10635_ _10636_ sky130_fd_sc_hd__o22a_2
X_12384_ VGND VPWR enc_block.round_key\[24\] _07962_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_129_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_806 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_209_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1312 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14123_ VPWR VGND VGND VPWR _09474_ _09594_ _09348_ sky130_fd_sc_hd__nor2_2
XFILLER_0_50_766 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19980_ VGND VPWR VPWR VGND _05400_ _11099_ keymem.key_mem\[10\]\[14\] _05406_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_183_2_Left_654 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_127_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18931_ VPWR VGND VGND VPWR _04654_ _04769_ _04179_ sky130_fd_sc_hd__nor2_2
XFILLER_0_265_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14054_ VGND VPWR VGND VPWR _09505_ _09429_ keymem.prev_key1_reg\[96\] _09526_ sky130_fd_sc_hd__a21o_2
X_13005_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[84\] _07843_ keymem.key_mem\[6\]\[84\]
+ _07639_ _08524_ sky130_fd_sc_hd__a22o_2
X_18862_ VPWR VGND _04707_ _04706_ enc_block.round_key\[43\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_20_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17813_ VGND VPWR _03187_ _09528_ _03804_ _03789_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_234_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18793_ VGND VPWR VPWR VGND _04600_ enc_block.block_w2_reg\[4\] _04030_ _04645_ sky130_fd_sc_hd__mux2_2
XFILLER_0_118_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17744_ VGND VPWR _00179_ _03760_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_222_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14956_ enc_block.sword_ctr_reg\[1\] _10420_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[13\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_262_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_76_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13907_ VPWR VGND VPWR VGND _09280_ _09291_ _09285_ _09338_ _09379_ sky130_fd_sc_hd__or4_2
XFILLER_0_37_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17675_ VGND VPWR VPWR VGND _03691_ key[145] keymem.prev_key1_reg\[17\] _03713_ sky130_fd_sc_hd__mux2_2
XFILLER_0_216_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14887_ VPWR VGND VPWR VGND _09664_ _10351_ _10352_ _09179_ _10350_ sky130_fd_sc_hd__or4b_2
XFILLER_0_37_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19414_ VGND VPWR VGND VPWR _05103_ keymem.key_mem_we _10284_ _05093_ _00506_ sky130_fd_sc_hd__a31o_2
X_16626_ VGND VPWR VGND VPWR _02780_ _02779_ _02782_ _02781_ sky130_fd_sc_hd__a21oi_2
X_13838_ VPWR VGND VPWR VGND _09307_ _09309_ _09285_ _09306_ _09310_ sky130_fd_sc_hd__or4_2
XFILLER_0_216_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19345_ VGND VPWR _00483_ _05057_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16557_ VGND VPWR VGND VPWR _02713_ _02712_ _02716_ _02714_ sky130_fd_sc_hd__a21oi_2
X_13769_ enc_block.sword_ctr_reg\[1\] _09241_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[24\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_45_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15508_ VGND VPWR _10968_ keymem.prev_key1_reg\[108\] _10917_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_19276_ VGND VPWR VGND VPWR _05012_ keymem.key_mem_we _03393_ _04999_ _00459_ sky130_fd_sc_hd__a31o_2
XFILLER_0_57_398 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16488_ VGND VPWR VGND VPWR _02649_ _09931_ _09796_ key[23] sky130_fd_sc_hd__o21a_2
X_18227_ VGND VPWR VGND VPWR _04135_ _04004_ _11089_ _11072_ sky130_fd_sc_hd__o21a_2
X_15439_ VPWR VGND VPWR VGND _10900_ key[11] _08936_ sky130_fd_sc_hd__or2_2
XFILLER_0_26_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18158_ VPWR VGND _04072_ _04071_ enc_block.round_key\[104\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_108_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_744 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_223_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17109_ VPWR VGND VGND VPWR _03225_ key[196] _08930_ sky130_fd_sc_hd__nand2_2
X_18089_ VGND VPWR _04008_ _03981_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_1_830 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_68_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_276 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20120_ VGND VPWR VPWR VGND _05469_ _03339_ keymem.key_mem\[10\]\[81\] _05479_ sky130_fd_sc_hd__mux2_2
XFILLER_0_110_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_141_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_885 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_1242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_81_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20051_ VGND VPWR VPWR VGND _05435_ _03035_ keymem.key_mem\[10\]\[48\] _05443_ sky130_fd_sc_hd__mux2_2
XFILLER_0_42_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23810_ VGND VPWR VPWR VGND clk _00303_ reset_n enc_block.block_w0_reg\[29\] sky130_fd_sc_hd__dfrtp_2
X_24790_ VGND VPWR VPWR VGND clk _01283_ reset_n keymem.key_mem\[6\]\[15\] sky130_fd_sc_hd__dfrtp_2
X_23741_ keymem.prev_key0_reg\[97\] clk _00238_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20953_ VGND VPWR _01225_ _05923_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_36_1013 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20884_ VPWR VGND keymem.key_mem\[7\]\[53\] _05887_ _05886_ VPWR VGND sky130_fd_sc_hd__and2_2
X_23672_ keymem.prev_key0_reg\[28\] clk _00169_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_88_1_Right_689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_48_321 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_220_271 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25411_ VGND VPWR VPWR VGND clk _01904_ reset_n keymem.key_mem\[2\]\[124\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_113_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22623_ VGND VPWR _02037_ _06781_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_48_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_165_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_516 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22554_ VGND VPWR _01987_ _06762_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25342_ VGND VPWR VPWR VGND clk _01835_ reset_n keymem.key_mem\[2\]\[55\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_48_398 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_118_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21505_ VGND VPWR _01485_ _06215_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_763 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22485_ VGND VPWR _01945_ _06735_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25273_ VGND VPWR VPWR VGND clk _01766_ reset_n keymem.key_mem\[3\]\[114\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_210_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_17_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24224_ VGND VPWR VPWR VGND clk _00717_ reset_n keymem.key_mem\[11\]\[89\] sky130_fd_sc_hd__dfrtp_2
X_21436_ VGND VPWR _01452_ _06179_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_228_1367 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_133_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24155_ VGND VPWR VPWR VGND clk _00648_ reset_n keymem.key_mem\[11\]\[20\] sky130_fd_sc_hd__dfrtp_2
X_21367_ VGND VPWR _01419_ _06143_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_31_265 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20318_ VGND VPWR VPWR VGND _05580_ _03006_ keymem.key_mem\[9\]\[45\] _05585_ sky130_fd_sc_hd__mux2_2
X_23106_ VGND VPWR VGND VPWR _02271_ _07030_ _07010_ keymem.prev_key1_reg\[94\] sky130_fd_sc_hd__o21a_2
X_24086_ VGND VPWR VPWR VGND clk _00579_ reset_n keymem.key_mem\[12\]\[79\] sky130_fd_sc_hd__dfrtp_2
X_21298_ VGND VPWR _01388_ _06105_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_120_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23037_ VGND VPWR VPWR VGND _06960_ _06988_ keymem.prev_key1_reg\[67\] _06989_ sky130_fd_sc_hd__mux2_2
XFILLER_0_124_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20249_ VGND VPWR VPWR VGND _05546_ _10977_ keymem.key_mem\[9\]\[12\] _05549_ sky130_fd_sc_hd__mux2_2
XFILLER_0_21_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_200_1242 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_198_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14810_ VGND VPWR VPWR VGND _10276_ keymem.prev_key1_reg\[70\] _10273_ _10274_ _09729_
+ sky130_fd_sc_hd__o31a_2
X_15790_ VGND VPWR _11246_ _11245_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24988_ VGND VPWR VPWR VGND clk _01481_ reset_n keymem.key_mem\[5\]\[85\] sky130_fd_sc_hd__dfrtp_2
X_14741_ VGND VPWR VGND VPWR _09132_ _09053_ _09687_ _09125_ _10207_ sky130_fd_sc_hd__o22a_2
X_23939_ VGND VPWR VPWR VGND clk _00432_ reset_n keymem.key_mem\[13\]\[60\] sky130_fd_sc_hd__dfrtp_2
X_11953_ VGND VPWR _07556_ _07555_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_19_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_265 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_233_1040 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17460_ VGND VPWR VGND VPWR _03282_ _02342_ _03537_ _03536_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_196_440 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14672_ VPWR VGND VPWR VGND _09768_ _10138_ _10139_ _09438_ _09446_ sky130_fd_sc_hd__or4b_2
XFILLER_0_98_298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_131_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_197_974 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11884_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[13\] dec_new_block\[109\]
+ _07506_ sky130_fd_sc_hd__mux2_2
XFILLER_0_170_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16411_ VPWR VGND VPWR VGND _02379_ _02523_ _02381_ _02378_ _02573_ sky130_fd_sc_hd__or4_2
X_13623_ VGND VPWR _09095_ _09094_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25609_ VGND VPWR VPWR VGND clk _02102_ reset_n keymem.key_mem\[0\]\[66\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_200_956 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17391_ VGND VPWR VGND VPWR _03477_ _03476_ _09791_ _10278_ sky130_fd_sc_hd__o21a_2
XFILLER_0_131_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19130_ VGND VPWR _00404_ _04921_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16342_ VGND VPWR VGND VPWR _11420_ _11296_ _11404_ _02505_ sky130_fd_sc_hd__a21o_2
X_13554_ VPWR VGND VPWR VGND _09026_ enc_block.block_w0_reg\[0\] _08952_ sky130_fd_sc_hd__or2_2
XFILLER_0_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12505_ VPWR VGND VPWR VGND _08072_ keymem.key_mem\[10\]\[35\] _07876_ keymem.key_mem\[12\]\[35\]
+ _07894_ _08073_ sky130_fd_sc_hd__a221o_2
X_19061_ VPWR VGND keymem.key_mem\[13\]\[2\] _04883_ _04880_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16273_ VPWR VGND VGND VPWR _11379_ _02437_ _11250_ sky130_fd_sc_hd__nor2_2
XFILLER_0_42_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13485_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[2\] _08956_ _08957_ _08943_ _08950_
+ _08953_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_120_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18012_ VPWR VGND VPWR VGND _03940_ _03729_ _03939_ sky130_fd_sc_hd__or2_2
X_15224_ VGND VPWR VGND VPWR _10686_ _10685_ _10687_ _10684_ _10683_ sky130_fd_sc_hd__nand4_2
XFILLER_0_168_1292 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_63_891 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12436_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[29\] _07668_ keymem.key_mem\[3\]\[29\]
+ _08009_ _08010_ sky130_fd_sc_hd__a22o_2
XFILLER_0_164_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15155_ VPWR VGND VGND VPWR _10619_ _10440_ _10477_ sky130_fd_sc_hd__nand2_2
X_12367_ VPWR VGND VPWR VGND _07946_ keymem.key_mem\[7\]\[23\] _07702_ keymem.key_mem\[9\]\[23\]
+ _07918_ _07947_ sky130_fd_sc_hd__a221o_2
XFILLER_0_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14106_ VGND VPWR VGND VPWR _09294_ _09396_ _09363_ _09311_ _09373_ _09577_ sky130_fd_sc_hd__o32a_2
XFILLER_0_61_1139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_142_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15086_ VPWR VGND VPWR VGND _10550_ _10474_ _10475_ _10541_ _10548_ _10549_ sky130_fd_sc_hd__o311a_2
X_12298_ VGND VPWR enc_block.round_key\[17\] _07883_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19963_ VGND VPWR _00762_ _05396_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_142_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18914_ VPWR VGND _04753_ enc_block.block_w3_reg\[23\] enc_block.block_w3_reg\[16\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_14037_ VGND VPWR VGND VPWR _09508_ _08932_ _09509_ _08937_ sky130_fd_sc_hd__nand3_2
XFILLER_0_266_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_129_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_105 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19894_ VGND VPWR _00731_ _05358_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_235_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18845_ VGND VPWR _04691_ _04086_ _00349_ _04602_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_101_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_886 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_173_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18776_ VPWR VGND VPWR VGND _04629_ _04625_ _04628_ sky130_fd_sc_hd__or2_2
XFILLER_0_235_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15988_ VGND VPWR VGND VPWR _11443_ _10732_ _11161_ _11441_ _11444_ sky130_fd_sc_hd__a31o_2
XFILLER_0_253_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17727_ VGND VPWR VGND VPWR _03732_ keymem.prev_key1_reg\[31\] _03751_ _03733_ sky130_fd_sc_hd__a21oi_2
X_14939_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[10\] _10402_ _10403_ _09255_ _10400_
+ _10401_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_54_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17658_ VGND VPWR _00152_ _03701_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_159_142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_153_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16609_ VGND VPWR VPWR VGND _02662_ keymem.key_mem\[14\]\[27\] _02765_ _02766_ sky130_fd_sc_hd__mux2_2
XFILLER_0_174_112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17589_ VGND VPWR _00136_ _03648_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_50_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19328_ VGND VPWR _05046_ _04876_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_50_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_2_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19259_ VPWR VGND keymem.key_mem_we _05002_ _03339_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_33_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_115_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_722 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22270_ VGND VPWR VPWR VGND _06622_ _03172_ keymem.key_mem\[2\]\[62\] _06624_ sky130_fd_sc_hd__mux2_2
XFILLER_0_260_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21221_ VGND VPWR _06065_ _05970_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_78_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_574 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_229_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21152_ VGND VPWR _06029_ _05971_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_160_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_660 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_121_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20103_ VGND VPWR _00828_ _05470_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_258_1305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21083_ VGND VPWR VPWR VGND _05983_ _02339_ keymem.key_mem\[6\]\[18\] _05993_ sky130_fd_sc_hd__mux2_2
XFILLER_0_0_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_499 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20034_ VGND VPWR VPWR VGND _05424_ _02955_ keymem.key_mem\[10\]\[40\] _05434_ sky130_fd_sc_hd__mux2_2
X_24911_ VGND VPWR VPWR VGND clk _01404_ reset_n keymem.key_mem\[5\]\[8\] sky130_fd_sc_hd__dfrtp_2
X_24842_ VGND VPWR VPWR VGND clk _01335_ reset_n keymem.key_mem\[6\]\[67\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24773_ VGND VPWR VPWR VGND clk _01266_ reset_n keymem.key_mem\[7\]\[126\] sky130_fd_sc_hd__dfrtp_2
X_21985_ VGND VPWR VGND VPWR _06472_ keymem.key_mem_we _03109_ _06446_ _01708_ sky130_fd_sc_hd__a31o_2
XFILLER_0_200_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23724_ keymem.prev_key0_reg\[80\] clk _00221_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20936_ VGND VPWR _01217_ _05914_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_138_326 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23655_ keymem.prev_key0_reg\[11\] clk _00152_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20867_ VGND VPWR _01185_ _05877_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_1141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22606_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[116\] _06777_ _06776_ _05066_ _02024_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_36_324 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23586_ VGND VPWR VPWR VGND clk _00087_ reset_n keymem.key_mem\[14\]\[75\] sky130_fd_sc_hd__dfrtp_2
X_20798_ VGND VPWR VGND VPWR _05840_ keymem.key_mem_we _11040_ _05838_ _01153_ sky130_fd_sc_hd__a31o_2
XFILLER_0_187_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_793 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25325_ VGND VPWR VPWR VGND clk _01818_ reset_n keymem.key_mem\[2\]\[38\] sky130_fd_sc_hd__dfrtp_2
X_22537_ VPWR VGND VGND VPWR _06757_ keymem.key_mem\[1\]\[68\] _06756_ sky130_fd_sc_hd__nand2_2
XFILLER_0_10_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_392 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_106_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25256_ VGND VPWR VPWR VGND clk _01749_ reset_n keymem.key_mem\[3\]\[97\] sky130_fd_sc_hd__dfrtp_2
X_13270_ VPWR VGND VPWR VGND _08762_ keymem.key_mem\[10\]\[110\] _07629_ keymem.key_mem\[1\]\[110\]
+ _07800_ _08763_ sky130_fd_sc_hd__a221o_2
X_22468_ VGND VPWR _01935_ _06728_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_106_289 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24207_ VGND VPWR VPWR VGND clk _00700_ reset_n keymem.key_mem\[11\]\[72\] sky130_fd_sc_hd__dfrtp_2
X_12221_ VGND VPWR _07812_ _07586_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21419_ VGND VPWR _01444_ _06170_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25187_ VGND VPWR VPWR VGND clk _01680_ reset_n keymem.key_mem\[3\]\[28\] sky130_fd_sc_hd__dfrtp_2
X_22399_ VGND VPWR VPWR VGND _06553_ _03647_ keymem.key_mem\[2\]\[124\] _06691_ sky130_fd_sc_hd__mux2_2
X_12152_ VGND VPWR _07748_ _07568_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24138_ VGND VPWR VPWR VGND clk _00631_ reset_n keymem.key_mem\[11\]\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_249_967 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16960_ VGND VPWR VGND VPWR _08930_ key[182] _03089_ _03090_ sky130_fd_sc_hd__a21o_2
X_12083_ VGND VPWR VGND VPWR _07600_ keymem.key_mem\[11\]\[4\] _07679_ _07681_ _07682_
+ _07572_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_21_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24069_ VGND VPWR VPWR VGND clk _00562_ reset_n keymem.key_mem\[12\]\[62\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_263_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_236_639 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15911_ VGND VPWR _11367_ _11361_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_229_691 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_21_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16891_ VGND VPWR _03027_ _09543_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_263_458 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_217_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_200_1061 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18630_ VGND VPWR _04498_ _04427_ _04435_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15842_ VGND VPWR _11298_ _11297_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_95_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_204_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_95_1279 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_176_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18561_ VGND VPWR _04436_ enc_block.block_w0_reg\[5\] _04435_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15773_ VGND VPWR _11229_ _11202_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12985_ VPWR VGND VPWR VGND _08505_ keymem.key_mem\[11\]\[82\] _07912_ keymem.key_mem\[1\]\[82\]
+ _07737_ _08506_ sky130_fd_sc_hd__a221o_2
XFILLER_0_8_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17512_ VGND VPWR _00126_ _03581_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14724_ VGND VPWR VPWR VGND _10190_ _10191_ _10189_ _10147_ _10187_ sky130_fd_sc_hd__a31oi_2
X_18492_ VGND VPWR _04374_ enc_block.block_w1_reg\[30\] _04373_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_11936_ VGND VPWR _07539_ _07538_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_59_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_262_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17443_ VPWR VGND VPWR VGND _03522_ _10737_ _10738_ sky130_fd_sc_hd__or2_2
X_14655_ VPWR VGND VGND VPWR _09749_ _10122_ _09401_ sky130_fd_sc_hd__nor2_2
XFILLER_0_135_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11867_ VGND VPWR result[100] _07497_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_129_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13606_ VPWR VGND VGND VPWR _09069_ _09078_ _09077_ sky130_fd_sc_hd__nor2_2
X_17374_ VGND VPWR VPWR VGND _03029_ _09508_ key[96] _03462_ sky130_fd_sc_hd__mux2_2
X_14586_ VGND VPWR VGND VPWR _09456_ _09302_ _09401_ _09426_ _09368_ _10054_ sky130_fd_sc_hd__o32a_2
XFILLER_0_39_184 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11798_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[2\] dec_new_block\[66\]
+ _07463_ sky130_fd_sc_hd__mux2_2
XFILLER_0_6_218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_54_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_131_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19113_ VPWR VGND keymem.key_mem\[13\]\[25\] _04912_ _04903_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_32_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16325_ _02486_ _02488_ _02484_ _02487_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_13537_ VGND VPWR _09009_ _09008_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_54_165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19044_ VGND VPWR _04869_ enc_block.block_w3_reg\[22\] _04868_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_16256_ VGND VPWR VGND VPWR _02420_ _11390_ _11389_ _11595_ _11491_ sky130_fd_sc_hd__a211o_2
X_13468_ VGND VPWR _08940_ _08939_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_67_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15207_ VGND VPWR VGND VPWR _10635_ _10668_ _10508_ _10563_ _10562_ _10670_ sky130_fd_sc_hd__o32a_2
XFILLER_0_112_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_208 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12419_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[28\] _07799_ keymem.key_mem\[2\]\[28\]
+ _07732_ _07994_ sky130_fd_sc_hd__a22o_2
XFILLER_0_2_435 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16187_ VGND VPWR VGND VPWR _02352_ _11323_ _11611_ _11355_ sky130_fd_sc_hd__o21a_2
XFILLER_0_51_872 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13399_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[123\] _07602_ keymem.key_mem\[7\]\[123\]
+ _07567_ _08879_ sky130_fd_sc_hd__a22o_2
X_15138_ VGND VPWR _10602_ _10601_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_142_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_241 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_120_270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15069_ VPWR VGND VPWR VGND _10505_ _10532_ _10512_ _10499_ _10533_ sky130_fd_sc_hd__or4_2
XFILLER_0_103_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19946_ VPWR VGND _05240_ _05386_ _05385_ VPWR VGND sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_178_1_Left_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_142_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_146_2_Left_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_103_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19877_ VGND VPWR _00723_ _05349_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_177_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18828_ VPWR VGND VGND VPWR _04676_ _04603_ _04675_ sky130_fd_sc_hd__nand2_2
XFILLER_0_78_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_218_1355 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18759_ VPWR VGND VGND VPWR _04613_ _04614_ _03994_ sky130_fd_sc_hd__nor2_2
XFILLER_0_77_202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21770_ VGND VPWR VPWR VGND _06355_ _03383_ keymem.key_mem\[4\]\[86\] _06356_ sky130_fd_sc_hd__mux2_2
XFILLER_0_81_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20721_ VGND VPWR VPWR VGND _05794_ _03543_ keymem.key_mem\[8\]\[108\] _05797_ sky130_fd_sc_hd__mux2_2
XFILLER_0_153_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23440_ VGND VPWR _07307_ _07085_ _07306_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20652_ VGND VPWR VGND VPWR _05676_ _03287_ _01087_ _05760_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_188_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_110_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_806 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23371_ VGND VPWR _07245_ _04159_ _02321_ _07096_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_50_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20583_ VGND VPWR _01054_ _05724_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_2_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_85_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25110_ VGND VPWR VPWR VGND clk _01603_ reset_n keymem.key_mem\[4\]\[79\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22322_ VGND VPWR VPWR VGND _06647_ _03392_ keymem.key_mem\[2\]\[87\] _06651_ sky130_fd_sc_hd__mux2_2
XFILLER_0_264_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_80 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1162 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22253_ VGND VPWR VPWR VGND _06611_ _03090_ keymem.key_mem\[2\]\[54\] _06615_ sky130_fd_sc_hd__mux2_2
X_25041_ VGND VPWR VPWR VGND clk _01534_ reset_n keymem.key_mem\[4\]\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_264_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_108_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21204_ VGND VPWR _06056_ _03287_ _01343_ _05985_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_22184_ VGND VPWR VPWR VGND _06578_ _02549_ keymem.key_mem\[2\]\[21\] _06579_ sky130_fd_sc_hd__mux2_2
XFILLER_0_125_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_160_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_252 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21135_ VGND VPWR _01310_ _06020_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_78_2_Left_549 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_111_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_121_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_160_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21066_ VGND VPWR VPWR VGND _05983_ _10835_ keymem.key_mem\[6\]\[10\] _05984_ sky130_fd_sc_hd__mux2_2
XFILLER_0_22_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_801 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20017_ VGND VPWR _00787_ _05425_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_96_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24825_ VGND VPWR VPWR VGND clk _01318_ reset_n keymem.key_mem\[6\]\[50\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_214_878 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_236_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_224 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12770_ VGND VPWR VGND VPWR _08313_ _07712_ keymem.key_mem\[6\]\[60\] _08310_ _08312_
+ sky130_fd_sc_hd__a211o_2
X_24756_ VGND VPWR VPWR VGND clk _01249_ reset_n keymem.key_mem\[7\]\[109\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_68_235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21968_ VGND VPWR _01700_ _06463_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_68_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11721_ VGND VPWR result[27] _07424_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_132_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23707_ keymem.prev_key0_reg\[63\] clk _00204_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20919_ VGND VPWR VGND VPWR _05905_ keymem.key_mem_we _03235_ _05893_ _01209_ sky130_fd_sc_hd__a31o_2
XFILLER_0_230_1032 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_192_2_Left_663 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_171_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24687_ VGND VPWR VPWR VGND clk _01180_ reset_n keymem.key_mem\[7\]\[40\] sky130_fd_sc_hd__dfrtp_2
X_21899_ VPWR VGND keymem.key_mem\[3\]\[17\] _06426_ _06413_ VPWR VGND sky130_fd_sc_hd__and2_2
X_14440_ VPWR VGND VPWR VGND _09904_ _09908_ _09909_ _09899_ _09902_ sky130_fd_sc_hd__or4b_2
XFILLER_0_132_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23638_ VGND VPWR VPWR VGND clk _00139_ reset_n keymem.key_mem\[14\]\[127\] sky130_fd_sc_hd__dfrtp_2
X_11652_ VGND VPWR VGND VPWR _07388_ keymem.round_ctr_reg\[3\] _07389_ keymem.round_ctr_reg\[1\]
+ _07387_ sky130_fd_sc_hd__nand4_2
XFILLER_0_167_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14371_ VPWR VGND VGND VPWR _09114_ _09204_ _09841_ _09658_ _09103_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_24_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23569_ VGND VPWR VPWR VGND clk _00070_ reset_n keymem.key_mem\[14\]\[58\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_153_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16110_ VGND VPWR VGND VPWR _11564_ _11222_ _11395_ _11266_ _11167_ sky130_fd_sc_hd__and4_2
XFILLER_0_153_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_51_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13322_ VPWR VGND VPWR VGND _08809_ keymem.key_mem\[3\]\[115\] _07690_ keymem.key_mem\[2\]\[115\]
+ _07647_ _08810_ sky130_fd_sc_hd__a221o_2
X_25308_ VGND VPWR VPWR VGND clk _01801_ reset_n keymem.key_mem\[2\]\[21\] sky130_fd_sc_hd__dfrtp_2
X_17090_ VPWR VGND VGND VPWR _03205_ _03206_ _03207_ _02866_ _03208_ sky130_fd_sc_hd__and4b_2
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16041_ VPWR VGND VPWR VGND _11495_ _11496_ _11493_ _11494_ sky130_fd_sc_hd__or3b_2
XFILLER_0_51_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_243_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25239_ VGND VPWR VPWR VGND clk _01732_ reset_n keymem.key_mem\[3\]\[80\] sky130_fd_sc_hd__dfrtp_2
X_13253_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[108\] _07565_ keymem.key_mem\[12\]\[108\]
+ _07787_ _08748_ sky130_fd_sc_hd__a22o_2
XFILLER_0_161_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12204_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[11\] _07577_ keymem.key_mem\[2\]\[11\]
+ _07545_ _07796_ sky130_fd_sc_hd__a22o_2
XFILLER_0_62_1234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13184_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[101\] _08577_ _08685_ _08681_ _08686_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_248_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_143_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19800_ VGND VPWR _00686_ _05309_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_209_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12135_ VGND VPWR _07731_ _07730_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_202_1134 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_202_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17992_ VGND VPWR VGND VPWR _03736_ keymem.prev_key0_reg\[120\] _03926_ _00261_ sky130_fd_sc_hd__a21o_2
XFILLER_0_40_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16943_ VPWR VGND VPWR VGND _03074_ _03071_ _03070_ key[180] _03027_ _03075_ sky130_fd_sc_hd__a221o_2
XFILLER_0_100_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19731_ VGND VPWR _00653_ _05273_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12066_ VGND VPWR _07666_ _07583_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_264_767 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1093 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16874_ VGND VPWR VGND VPWR _11051_ _11050_ _03012_ _03011_ sky130_fd_sc_hd__a21oi_2
X_19662_ VGND VPWR VPWR VGND _05227_ _05081_ keymem.key_mem\[12\]\[123\] _05235_ sky130_fd_sc_hd__mux2_2
XFILLER_0_204_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_232_620 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_126_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_254_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15825_ VPWR VGND VPWR VGND _11264_ _11216_ _11179_ _11232_ _11281_ sky130_fd_sc_hd__or4_2
X_18613_ VPWR VGND VGND VPWR _04482_ _04483_ _04478_ sky130_fd_sc_hd__nor2_2
XFILLER_0_260_951 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19593_ VPWR VGND keymem.key_mem\[12\]\[90\] _05199_ _05173_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_204_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15756_ enc_block.sword_ctr_reg\[1\] _11212_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[16\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_18544_ VPWR VGND VPWR VGND _04420_ block[75] _04330_ enc_block.block_w3_reg\[11\]
+ _04276_ _04421_ sky130_fd_sc_hd__a221o_2
XFILLER_0_99_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12968_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[80\] _07683_ keymem.key_mem\[3\]\[80\]
+ _07603_ _08491_ sky130_fd_sc_hd__a22o_2
XFILLER_0_220_848 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_231_196 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14707_ VPWR VGND VGND VPWR _09100_ _10174_ _09136_ sky130_fd_sc_hd__nor2_2
XFILLER_0_59_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11919_ VGND VPWR result[126] _07523_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18475_ _04357_ _04359_ _04065_ _04358_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_206_91 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_169_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_150_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15687_ VGND VPWR _11144_ keymem.prev_key0_reg\[111\] _11143_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_12899_ VGND VPWR VGND VPWR _07584_ keymem.key_mem\[14\]\[73\] _08425_ _08427_ _08429_
+ _08428_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_111_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17426_ VGND VPWR _00114_ _03507_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14638_ VGND VPWR VGND VPWR _09333_ _09565_ _09341_ _09419_ _10105_ sky130_fd_sc_hd__o22a_2
XFILLER_0_150_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_111_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17357_ VGND VPWR VGND VPWR _02822_ _02817_ _03447_ _03446_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_144_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14569_ VGND VPWR VGND VPWR _09378_ _09415_ _09330_ _09749_ _10037_ sky130_fd_sc_hd__o22a_2
XFILLER_0_248_1359 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16308_ VPWR VGND VPWR VGND _02472_ keymem.prev_key1_reg\[84\] sky130_fd_sc_hd__inv_2
XFILLER_0_27_198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17288_ VGND VPWR _00098_ _03385_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_67_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_43_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19027_ VGND VPWR _04854_ enc_block.block_w3_reg\[21\] enc_block.block_w1_reg\[5\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16239_ VGND VPWR _09729_ keymem.prev_key1_reg\[19\] _02404_ keymem.prev_key1_reg\[51\]
+ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_261_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_321 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_2_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_152_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_23_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_267_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_76_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19929_ VGND VPWR VPWR VGND _05372_ keymem.key_mem\[11\]\[120\] _03620_ _05377_ sky130_fd_sc_hd__mux2_2
XFILLER_0_208_650 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_76_96 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22940_ VGND VPWR VPWR VGND _06914_ _06931_ keymem.prev_key1_reg\[27\] _06932_ sky130_fd_sc_hd__mux2_2
XFILLER_0_78_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_190_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22871_ VGND VPWR VGND VPWR _09929_ _03795_ _06887_ _09990_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_39_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24610_ VGND VPWR VPWR VGND clk _01103_ reset_n keymem.key_mem\[8\]\[91\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_210_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21822_ VGND VPWR VPWR VGND _06377_ _03560_ keymem.key_mem\[4\]\[111\] _06383_ sky130_fd_sc_hd__mux2_2
X_25590_ VGND VPWR VPWR VGND clk _02083_ reset_n keymem.key_mem\[0\]\[47\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_210_336 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24541_ VGND VPWR VPWR VGND clk _01034_ reset_n keymem.key_mem\[8\]\[22\] sky130_fd_sc_hd__dfrtp_2
X_21753_ VGND VPWR VPWR VGND _06344_ _03314_ keymem.key_mem\[4\]\[78\] _06347_ sky130_fd_sc_hd__mux2_2
XFILLER_0_175_240 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20704_ VGND VPWR VPWR VGND _05783_ _03492_ keymem.key_mem\[8\]\[100\] _05788_ sky130_fd_sc_hd__mux2_2
X_24472_ VGND VPWR VPWR VGND clk _00965_ reset_n keymem.key_mem\[9\]\[81\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_18_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_46_430 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_114_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21684_ VGND VPWR VPWR VGND _06308_ _03006_ keymem.key_mem\[4\]\[45\] _06311_ sky130_fd_sc_hd__mux2_2
X_23423_ VGND VPWR _07292_ _07231_ _07291_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20635_ VGND VPWR VPWR VGND _05747_ _03216_ keymem.key_mem\[8\]\[67\] _05752_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_34_614 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_149_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23354_ VGND VPWR VGND VPWR _07230_ _03992_ _07228_ _07229_ _02319_ sky130_fd_sc_hd__a31o_2
XFILLER_0_116_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20566_ VGND VPWR VPWR VGND _05714_ _02893_ keymem.key_mem\[8\]\[34\] _05716_ sky130_fd_sc_hd__mux2_2
XFILLER_0_190_276 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_149_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_85_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22305_ VGND VPWR VPWR VGND _06634_ _03321_ keymem.key_mem\[2\]\[79\] _06642_ sky130_fd_sc_hd__mux2_2
X_23285_ VGND VPWR _07168_ enc_block.block_w0_reg\[16\] _07167_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20497_ VGND VPWR _05679_ _05675_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_371 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25024_ VGND VPWR VPWR VGND clk _01517_ reset_n keymem.key_mem\[5\]\[121\] sky130_fd_sc_hd__dfrtp_2
X_22236_ VGND VPWR VPWR VGND _06600_ _03015_ keymem.key_mem\[2\]\[46\] _06606_ sky130_fd_sc_hd__mux2_2
XFILLER_0_221_1009 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_203_1410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22167_ VGND VPWR VPWR VGND _06565_ _11039_ keymem.key_mem\[2\]\[13\] _06570_ sky130_fd_sc_hd__mux2_2
X_21118_ VGND VPWR _01302_ _06011_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22098_ VGND VPWR VPWR VGND _06527_ _05054_ keymem.key_mem\[3\]\[110\] _06532_ sky130_fd_sc_hd__mux2_2
XFILLER_0_22_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13940_ VGND VPWR VGND VPWR _09336_ _09386_ _09411_ _09408_ _09412_ sky130_fd_sc_hd__o22a_2
X_21049_ VGND VPWR VPWR VGND _05972_ _09861_ keymem.key_mem\[6\]\[2\] _05975_ sky130_fd_sc_hd__mux2_2
XFILLER_0_199_811 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_439 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_96_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13871_ VGND VPWR _09343_ _09342_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_9_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15610_ VPWR VGND VGND VPWR _11068_ _11066_ _11067_ sky130_fd_sc_hd__nand2_2
XFILLER_0_57_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12822_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[66\] _07748_ keymem.key_mem\[10\]\[66\]
+ _07876_ _08359_ sky130_fd_sc_hd__a22o_2
X_24808_ VGND VPWR VPWR VGND clk _01301_ reset_n keymem.key_mem\[6\]\[33\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_213_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16590_ VGND VPWR VGND VPWR _02393_ _02745_ _02747_ _02372_ sky130_fd_sc_hd__nand3_2
XFILLER_0_9_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25788_ keymem.prev_key1_reg\[104\] clk _02281_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_232_1138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_202_859 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15541_ VPWR VGND VGND VPWR _10559_ _11000_ _10509_ sky130_fd_sc_hd__nor2_2
XFILLER_0_9_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12753_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[59\] _07844_ keymem.key_mem\[2\]\[59\]
+ _07698_ _08297_ sky130_fd_sc_hd__a22o_2
X_24739_ VGND VPWR VPWR VGND clk _01232_ reset_n keymem.key_mem\[7\]\[92\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_56_216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11704_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[19\] dec_new_block\[19\]
+ _07416_ sky130_fd_sc_hd__mux2_2
X_18260_ VPWR VGND VGND VPWR _04165_ _04162_ _04163_ sky130_fd_sc_hd__nand2_2
X_15472_ VPWR VGND VGND VPWR _10543_ _10639_ _10932_ _10867_ _10644_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_210_892 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12684_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[52\] _07668_ keymem.key_mem\[8\]\[52\]
+ _07878_ _08235_ sky130_fd_sc_hd__a22o_2
XFILLER_0_132_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17211_ VPWR VGND VGND VPWR _03316_ key[207] _10086_ sky130_fd_sc_hd__nand2_2
X_14423_ VGND VPWR VGND VPWR _09388_ _09391_ _09404_ _09381_ _09892_ sky130_fd_sc_hd__o22a_2
X_18191_ VPWR VGND VGND VPWR _04102_ _04098_ _04100_ sky130_fd_sc_hd__nand2_2
X_11635_ VGND VPWR VGND VPWR enc_block.enc_ctrl_reg\[0\] encdec _07375_ next sky130_fd_sc_hd__nand3_2
XFILLER_0_167_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17142_ VPWR VGND VPWR VGND _10379_ _10375_ key[200] _03077_ _03254_ sky130_fd_sc_hd__a22o_2
X_14354_ VGND VPWR VGND VPWR _09154_ _09221_ _09824_ _09178_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_68_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_128_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13305_ VGND VPWR enc_block.round_key\[113\] _08794_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_40_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17073_ VGND VPWR VGND VPWR _08930_ key[192] _03192_ _03193_ sky130_fd_sc_hd__a21o_2
X_14285_ VGND VPWR VGND VPWR _09426_ _09576_ _09754_ _09420_ _09755_ sky130_fd_sc_hd__o22a_2
XFILLER_0_29_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16024_ VGND VPWR VGND VPWR _11460_ _11420_ _11479_ _11379_ sky130_fd_sc_hd__a21oi_2
X_13236_ VGND VPWR enc_block.round_key\[106\] _08732_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_122_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_179_1_Right_780 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13167_ VPWR VGND VPWR VGND _08669_ keymem.key_mem\[5\]\[100\] _08096_ keymem.key_mem\[7\]\[100\]
+ _08050_ _08670_ sky130_fd_sc_hd__a221o_2
XFILLER_0_0_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_594 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12118_ VGND VPWR _07715_ _07714_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_178_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17975_ VGND VPWR VPWR VGND _03281_ key[243] keymem.prev_key1_reg\[115\] _03915_
+ sky130_fd_sc_hd__mux2_2
X_13098_ VPWR VGND VPWR VGND _08607_ keymem.key_mem\[9\]\[93\] _07717_ keymem.key_mem\[11\]\[93\]
+ _07781_ _08608_ sky130_fd_sc_hd__a221o_2
XFILLER_0_100_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19714_ VGND VPWR _00645_ _05264_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_139_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16926_ VPWR VGND VPWR VGND _03059_ _02399_ sky130_fd_sc_hd__inv_2
X_12049_ VGND VPWR _07649_ _07567_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_178_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_174_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_139_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19645_ VGND VPWR VPWR VGND _05216_ _05064_ keymem.key_mem\[12\]\[115\] _05226_ sky130_fd_sc_hd__mux2_2
XFILLER_0_79_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16857_ VPWR VGND VGND VPWR _02997_ key[172] _02875_ sky130_fd_sc_hd__nand2_2
XFILLER_0_75_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15808_ VGND VPWR VGND VPWR _11264_ _11171_ _11170_ keymem.prev_key1_reg\[19\] _08954_
+ _08941_ sky130_fd_sc_hd__a32o_2
X_16788_ VPWR VGND VPWR VGND _02933_ _02929_ _02926_ key[166] _02875_ _02934_ sky130_fd_sc_hd__a221o_2
X_19576_ VGND VPWR _00581_ _05190_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_1_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1194 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15739_ VGND VPWR VGND VPWR enc_block.block_w1_reg\[20\] _08985_ _10387_ _11193_
+ _11195_ _11194_ sky130_fd_sc_hd__a2111o_2
X_18527_ VPWR VGND _04406_ _04405_ enc_block.round_key\[73\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_48_728 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_62_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_47_216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18458_ VGND VPWR _04343_ enc_block.block_w0_reg\[2\] _04342_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17409_ VGND VPWR VPWR VGND _03467_ keymem.key_mem\[14\]\[100\] _03492_ _03493_ sky130_fd_sc_hd__mux2_2
XFILLER_0_8_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18389_ VPWR VGND _04282_ _04281_ enc_block.round_key\[125\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_111_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_271 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_185_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20420_ VGND VPWR _05638_ _05533_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_55_293 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_86_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_185_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20351_ VGND VPWR _05602_ _05533_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23070_ VGND VPWR VPWR VGND _06992_ _03328_ keymem.prev_key1_reg\[80\] _07009_ sky130_fd_sc_hd__mux2_2
XFILLER_0_113_376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20282_ VGND VPWR VPWR VGND _05558_ _02787_ keymem.key_mem\[9\]\[28\] _05566_ sky130_fd_sc_hd__mux2_2
XFILLER_0_144_1165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22021_ VGND VPWR VGND VPWR _06491_ keymem.key_mem_we _03268_ _06475_ _01725_ sky130_fd_sc_hd__a31o_2
XFILLER_0_122_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23972_ VGND VPWR VPWR VGND clk _00465_ reset_n keymem.key_mem\[13\]\[93\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25711_ keymem.prev_key1_reg\[27\] clk _02204_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_157_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22923_ VGND VPWR VPWR VGND _06914_ _06919_ keymem.prev_key1_reg\[22\] _06920_ sky130_fd_sc_hd__mux2_2
XFILLER_0_237_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25642_ VGND VPWR VPWR VGND clk _02135_ reset_n keymem.key_mem\[0\]\[99\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_233_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22854_ VGND VPWR _02174_ _06875_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_196_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1211 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_233_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21805_ VGND VPWR VPWR VGND _06366_ _03511_ keymem.key_mem\[4\]\[103\] _06374_ sky130_fd_sc_hd__mux2_2
XFILLER_0_6_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25573_ VGND VPWR VPWR VGND clk _02066_ reset_n keymem.key_mem\[0\]\[30\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22785_ VGND VPWR _02127_ _06853_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_151_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24524_ VGND VPWR VPWR VGND clk _01017_ reset_n keymem.key_mem\[8\]\[5\] sky130_fd_sc_hd__dfrtp_2
X_21736_ VGND VPWR VPWR VGND _06330_ _03245_ keymem.key_mem\[4\]\[70\] _06338_ sky130_fd_sc_hd__mux2_2
XFILLER_0_108_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_108_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24455_ VGND VPWR VPWR VGND clk _00948_ reset_n keymem.key_mem\[9\]\[64\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_163_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21667_ VGND VPWR VPWR VGND _06297_ _02923_ keymem.key_mem\[4\]\[37\] _06302_ sky130_fd_sc_hd__mux2_2
XFILLER_0_30_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23406_ VGND VPWR _07277_ _07204_ _07276_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20618_ VGND VPWR VPWR VGND _05736_ _03139_ keymem.key_mem\[8\]\[59\] _05743_ sky130_fd_sc_hd__mux2_2
XFILLER_0_62_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_227_1229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24386_ VGND VPWR VPWR VGND clk _00879_ reset_n keymem.key_mem\[10\]\[123\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_164_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_904 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21598_ VGND VPWR VPWR VGND _06263_ _10098_ keymem.key_mem\[4\]\[4\] _06266_ sky130_fd_sc_hd__mux2_2
XFILLER_0_123_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23337_ _07213_ _07215_ _07212_ _07214_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_61_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20549_ VGND VPWR VPWR VGND _05703_ _02742_ keymem.key_mem\[8\]\[26\] _05707_ sky130_fd_sc_hd__mux2_2
XFILLER_0_205_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14070_ VGND VPWR VPWR VGND _09541_ keymem.key_mem\[14\]\[0\] _09537_ _09542_ sky130_fd_sc_hd__mux2_2
X_23268_ _07151_ _07153_ _04103_ _07152_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_240_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_205_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13021_ VGND VPWR VGND VPWR _08539_ _07721_ keymem.key_mem\[14\]\[85\] _08536_ _08538_
+ sky130_fd_sc_hd__a211o_2
X_25007_ VGND VPWR VPWR VGND clk _01500_ reset_n keymem.key_mem\[5\]\[104\] sky130_fd_sc_hd__dfrtp_2
X_22219_ VGND VPWR VPWR VGND _06589_ _02934_ keymem.key_mem\[2\]\[38\] _06597_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_18_Left_286 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23199_ VPWR VGND VPWR VGND _07089_ block[0] _04351_ enc_block.block_w2_reg\[0\]
+ _03978_ _07090_ sky130_fd_sc_hd__a221o_2
XFILLER_0_246_520 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_918 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14972_ VPWR VGND VPWR VGND _10424_ _10435_ _10430_ _10419_ _10436_ sky130_fd_sc_hd__or4_2
X_17760_ VGND VPWR VPWR VGND _03763_ _03770_ keymem.prev_key0_reg\[44\] _03771_ sky130_fd_sc_hd__mux2_2
X_13923_ VPWR VGND VPWR VGND _09299_ _09246_ _09315_ _09297_ _09395_ sky130_fd_sc_hd__or4_2
X_16711_ VGND VPWR _00043_ _02863_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_96_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17691_ VGND VPWR VPWR VGND _03723_ _02604_ keymem.prev_key0_reg\[22\] _03724_ sky130_fd_sc_hd__mux2_2
XFILLER_0_57_1155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19430_ VPWR VGND keymem.key_mem\[12\]\[14\] _05112_ _05102_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16642_ VPWR VGND VPWR VGND _02797_ key[29] _09719_ sky130_fd_sc_hd__or2_2
XFILLER_0_18_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13854_ VPWR VGND VPWR VGND _09299_ _09245_ _09314_ _09254_ _09326_ sky130_fd_sc_hd__or4_2
XFILLER_0_251_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_198_162 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_212_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12805_ VPWR VGND VPWR VGND _08343_ keymem.key_mem\[5\]\[64\] _07780_ keymem.key_mem\[8\]\[64\]
+ _07753_ _08344_ sky130_fd_sc_hd__a221o_2
X_19361_ VGND VPWR _00488_ _05068_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16573_ VGND VPWR _02731_ _02728_ _02730_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_13785_ VGND VPWR VGND VPWR _09257_ enc_block.block_w2_reg\[26\] enc_block.sword_ctr_reg\[1\]
+ enc_block.sword_ctr_reg\[0\] sky130_fd_sc_hd__and3b_2
XPHY_EDGE_ROW_27_Left_295 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_241_Right_110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_186_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15524_ VPWR VGND VPWR VGND _10982_ _10983_ _10980_ _10770_ sky130_fd_sc_hd__or3b_2
X_18312_ VPWR VGND VPWR VGND _04212_ _04189_ _04210_ enc_block.block_w0_reg\[21\]
+ _04097_ _00295_ sky130_fd_sc_hd__a221o_2
XFILLER_0_96_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19292_ VGND VPWR VPWR VGND _04993_ _05021_ keymem.key_mem\[13\]\[94\] _05022_ sky130_fd_sc_hd__mux2_2
X_12736_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[57\] _07639_ keymem.key_mem\[10\]\[57\]
+ _08193_ _08282_ sky130_fd_sc_hd__a22o_2
XFILLER_0_29_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_267_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18243_ VGND VPWR VGND VPWR _04146_ enc_block.round_key\[111\] _04149_ _04150_ sky130_fd_sc_hd__a21o_2
XFILLER_0_38_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_187_1_Left_454 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15455_ VGND VPWR _10915_ keymem.prev_key0_reg\[44\] keymem.prev_key0_reg\[76\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
X_12667_ VGND VPWR VGND VPWR _08220_ _07665_ keymem.key_mem\[4\]\[50\] _08217_ _08219_
+ sky130_fd_sc_hd__a211o_2
X_14406_ VGND VPWR VGND VPWR _09875_ _09872_ _09871_ _09749_ _09874_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_245_1307 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_155_2_Left_626 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_742 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18174_ VPWR VGND VGND VPWR _04086_ _04087_ _04041_ sky130_fd_sc_hd__nor2_2
X_15386_ VPWR VGND VGND VPWR _10595_ _10847_ _10521_ sky130_fd_sc_hd__nor2_2
XFILLER_0_41_904 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_68_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12598_ VPWR VGND VPWR VGND _08156_ keymem.key_mem\[9\]\[44\] _07842_ keymem.key_mem\[10\]\[44\]
+ _07877_ _08157_ sky130_fd_sc_hd__a221o_2
XFILLER_0_29_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17125_ VGND VPWR VGND VPWR _10264_ _10263_ _03239_ _03237_ sky130_fd_sc_hd__a21oi_2
X_14337_ VPWR VGND VGND VPWR _09204_ _09168_ _09178_ _09153_ _09807_ _09806_ sky130_fd_sc_hd__o221a_2
XFILLER_0_53_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_499 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_52_285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17056_ VGND VPWR VPWR VGND _03175_ _02691_ _03177_ _09722_ _03176_ sky130_fd_sc_hd__o211a_2
X_14268_ VGND VPWR VGND VPWR _09737_ _09404_ _09419_ _09475_ _09738_ sky130_fd_sc_hd__a31o_2
XFILLER_0_21_650 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_204_1037 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16007_ VGND VPWR VGND VPWR _11236_ _11246_ _11400_ _11462_ sky130_fd_sc_hd__a21o_2
XFILLER_0_110_335 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13219_ VPWR VGND VPWR VGND _08716_ keymem.key_mem\[10\]\[105\] _07909_ keymem.key_mem\[4\]\[105\]
+ _07637_ _08717_ sky130_fd_sc_hd__a221o_2
X_14199_ _09190_ _09670_ _09181_ _09199_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_221_1340 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_104_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17958_ VGND VPWR _00250_ _03903_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_139_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16909_ VGND VPWR VGND VPWR _03041_ _03040_ _03043_ _03044_ sky130_fd_sc_hd__a21o_2
XFILLER_0_79_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17889_ VGND VPWR _00228_ _03856_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_75_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19628_ VGND VPWR _00606_ _05217_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_36_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19559_ VGND VPWR VPWR VGND _05151_ _04989_ keymem.key_mem\[12\]\[74\] _05181_ sky130_fd_sc_hd__mux2_2
XFILLER_0_215_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22570_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[89\] _06767_ _06766_ _05015_ _01997_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_8_622 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_2_Left_558 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21521_ VGND VPWR VPWR VGND _06220_ _03474_ keymem.key_mem\[5\]\[97\] _06224_ sky130_fd_sc_hd__mux2_2
XFILLER_0_56_580 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_267_1565 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_1248 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24240_ VGND VPWR VPWR VGND clk _00733_ reset_n keymem.key_mem\[11\]\[105\] sky130_fd_sc_hd__dfrtp_2
X_21452_ VGND VPWR VPWR VGND _06184_ _03193_ keymem.key_mem\[5\]\[64\] _06188_ sky130_fd_sc_hd__mux2_2
XFILLER_0_7_198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_298 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20403_ VGND VPWR _00969_ _05629_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_43_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21383_ VGND VPWR VPWR VGND _06151_ _02861_ keymem.key_mem\[5\]\[31\] _06152_ sky130_fd_sc_hd__mux2_2
X_24171_ VGND VPWR VPWR VGND clk _00664_ reset_n keymem.key_mem\[11\]\[36\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_850 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23122_ VGND VPWR _02277_ _07040_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20334_ VGND VPWR _00936_ _05593_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_113_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_101_324 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_970 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20265_ VGND VPWR VPWR VGND _05546_ _02480_ keymem.key_mem\[9\]\[20\] _05557_ sky130_fd_sc_hd__mux2_2
X_23053_ VGND VPWR VPWR VGND _06992_ _03266_ keymem.prev_key1_reg\[73\] _06999_ sky130_fd_sc_hd__mux2_2
X_22004_ VGND VPWR _01717_ _06482_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_200_1424 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_262_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20196_ VGND VPWR VPWR VGND _05515_ _03600_ keymem.key_mem\[10\]\[117\] _05519_ sky130_fd_sc_hd__mux2_2
XFILLER_0_157_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23955_ VGND VPWR VPWR VGND clk _00448_ reset_n keymem.key_mem\[13\]\[76\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_97_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_729 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_212_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22906_ VPWR VGND VPWR VGND _06909_ _11445_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23886_ VGND VPWR VPWR VGND clk _00379_ reset_n keymem.key_mem\[13\]\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25625_ VGND VPWR VPWR VGND clk _02118_ reset_n keymem.key_mem\[0\]\[82\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_233_1266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22837_ VGND VPWR VGND VPWR _02165_ _06866_ _06865_ keymem.rcon_logic.tmp_rcon\[2\]
+ _06867_ _06864_ sky130_fd_sc_hd__a32o_2
XFILLER_0_39_514 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_66_322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13570_ VPWR VGND VGND VPWR _09039_ _09042_ _09041_ sky130_fd_sc_hd__nor2_2
X_25556_ VGND VPWR VPWR VGND clk _02049_ reset_n keymem.key_mem\[0\]\[13\] sky130_fd_sc_hd__dfrtp_2
X_22768_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[81\] _06837_ _06836_ _05002_ _02117_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_136_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12521_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[37\] _07787_ keymem.key_mem\[4\]\[37\]
+ _07913_ _08087_ sky130_fd_sc_hd__a22o_2
X_24507_ VGND VPWR VPWR VGND clk _01000_ reset_n keymem.key_mem\[9\]\[116\] sky130_fd_sc_hd__dfrtp_2
X_21719_ VGND VPWR VPWR VGND _06319_ _03172_ keymem.key_mem\[4\]\[62\] _06329_ sky130_fd_sc_hd__mux2_2
XFILLER_0_66_388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25487_ VGND VPWR VPWR VGND clk _01980_ reset_n keymem.key_mem\[1\]\[72\] sky130_fd_sc_hd__dfrtp_2
X_22699_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[40\] _06790_ _06789_ _04935_ _02076_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_19_271 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15240_ VGND VPWR VPWR VGND _10478_ _10495_ _10514_ _10703_ sky130_fd_sc_hd__or3_2
XFILLER_0_129_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24438_ VGND VPWR VPWR VGND clk _00931_ reset_n keymem.key_mem\[9\]\[47\] sky130_fd_sc_hd__dfrtp_2
X_12452_ VGND VPWR VGND VPWR _08025_ _07580_ keymem.key_mem\[12\]\[30\] _08022_ _08024_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_168_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_213 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_191_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_50_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_69_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15171_ VGND VPWR _10635_ _10634_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_62_583 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12383_ VGND VPWR VGND VPWR _07793_ keymem.key_mem\[0\]\[24\] _07961_ _07956_ _07954_
+ _07962_ sky130_fd_sc_hd__o32a_2
X_24369_ VGND VPWR VPWR VGND clk _00862_ reset_n keymem.key_mem\[10\]\[106\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_65_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14122_ VGND VPWR VGND VPWR _09449_ _09357_ _09593_ _09329_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_209_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18930_ VPWR VGND _04768_ _04767_ enc_block.round_key\[50\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_127_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14053_ VGND VPWR _09524_ _09522_ _09525_ _09520_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_265_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13004_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[84\] _07650_ keymem.key_mem\[1\]\[84\]
+ _07901_ _08523_ sky130_fd_sc_hd__a22o_2
X_18861_ VPWR VGND VPWR VGND _04705_ block[43] _04576_ enc_block.block_w0_reg\[11\]
+ _04666_ _04706_ sky130_fd_sc_hd__a221o_2
XFILLER_0_94_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_101_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_197_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17812_ VPWR VGND VPWR VGND _03181_ _03803_ keymem.prev_key0_reg\[63\] _03788_ _00204_
+ sky130_fd_sc_hd__a22o_2
X_18792_ VPWR VGND _04644_ _04643_ enc_block.round_key\[36\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_175_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14955_ VGND VPWR VGND VPWR _10419_ _10418_ _10417_ keymem.prev_key1_reg\[12\] _10402_
+ _09255_ sky130_fd_sc_hd__a32o_2
XFILLER_0_76_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17743_ VGND VPWR VPWR VGND _03723_ _02931_ keymem.prev_key0_reg\[38\] _03760_ sky130_fd_sc_hd__mux2_2
XFILLER_0_136_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13906_ VGND VPWR _09378_ _09377_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_76_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_35_Left_303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14886_ VGND VPWR VGND VPWR _09080_ _09137_ _09077_ _09177_ _09040_ _10351_ sky130_fd_sc_hd__o32a_2
X_17674_ VGND VPWR _00157_ _03712_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_216_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19413_ VPWR VGND keymem.key_mem\[12\]\[6\] _05103_ _05102_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13837_ VGND VPWR _09309_ _09308_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_76_108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16625_ VPWR VGND _02781_ keymem.prev_key1_reg\[60\] keymem.prev_key1_reg\[28\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_251_1366 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_216_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19344_ VGND VPWR VPWR VGND _05046_ _05056_ keymem.key_mem\[13\]\[111\] _05057_ sky130_fd_sc_hd__mux2_2
X_16556_ _02713_ _02715_ _02712_ _02714_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_13768_ VGND VPWR _09240_ _07385_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_45_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15507_ VGND VPWR _10967_ _09522_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_112_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12719_ VPWR VGND VPWR VGND _08266_ keymem.key_mem\[13\]\[55\] _07730_ keymem.key_mem\[8\]\[55\]
+ _08265_ _08267_ sky130_fd_sc_hd__a221o_2
X_16487_ VGND VPWR _02647_ _02645_ _02648_ _02646_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_19275_ VPWR VGND keymem.key_mem\[13\]\[87\] _05012_ _04979_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_150_13 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13699_ VPWR VGND VPWR VGND _09045_ _09154_ _09015_ _09014_ _09171_ sky130_fd_sc_hd__or4_2
XFILLER_0_210_1074 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18226_ VPWR VGND VGND VPWR _04134_ enc_block.round_key\[110\] _04132_ sky130_fd_sc_hd__nand2_2
X_15438_ VGND VPWR VGND VPWR _10895_ _10894_ _10899_ _10897_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_216_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_186_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_775 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_147_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18157_ VPWR VGND VPWR VGND _04070_ block[104] _03959_ enc_block.block_w2_reg\[8\]
+ _03954_ _04071_ sky130_fd_sc_hd__a221o_2
X_15369_ VPWR VGND VGND VPWR _10831_ key[138] _10091_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_44_Left_312 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_83_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_222 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17108_ VGND VPWR VGND VPWR _03224_ _03222_ _02647_ _03223_ _10190_ sky130_fd_sc_hd__a211o_2
XFILLER_0_159_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18088_ VGND VPWR _04007_ _03977_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_29_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17039_ VGND VPWR _03162_ _03161_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_223_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1210 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_110_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20050_ VGND VPWR _00803_ _05442_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_258_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1254 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_256_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Left_321 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_84_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_154_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23740_ keymem.prev_key0_reg\[96\] clk _00237_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20952_ VGND VPWR VPWR VGND _05912_ _05008_ keymem.key_mem\[7\]\[85\] _05923_ sky130_fd_sc_hd__mux2_2
XFILLER_0_36_1025 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_234_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_812 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23671_ keymem.prev_key0_reg\[27\] clk _00168_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_152_1242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20883_ VGND VPWR _05886_ _05823_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25410_ VGND VPWR VPWR VGND clk _01903_ reset_n keymem.key_mem\[2\]\[123\] sky130_fd_sc_hd__dfrtp_2
X_22622_ VGND VPWR VPWR VGND _06779_ keymem.key_mem\[0\]\[1\] _09725_ _06781_ sky130_fd_sc_hd__mux2_2
XFILLER_0_165_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25341_ VGND VPWR VPWR VGND clk _01834_ reset_n keymem.key_mem\[2\]\[54\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_8_430 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22553_ VGND VPWR VPWR VGND _06750_ keymem.key_mem\[1\]\[79\] _03322_ _06762_ sky130_fd_sc_hd__mux2_2
XFILLER_0_1_1012 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21504_ VGND VPWR VPWR VGND _06209_ _03409_ keymem.key_mem\[5\]\[89\] _06215_ sky130_fd_sc_hd__mux2_2
X_25272_ VGND VPWR VPWR VGND clk _01765_ reset_n keymem.key_mem\[3\]\[113\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_1056 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_90_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_267_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22484_ VGND VPWR VPWR VGND _06726_ keymem.key_mem\[1\]\[37\] _02924_ _06735_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_62_Left_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_775 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_173_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_133_235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24223_ VGND VPWR VPWR VGND clk _00716_ reset_n keymem.key_mem\[11\]\[88\] sky130_fd_sc_hd__dfrtp_2
X_21435_ VGND VPWR VPWR VGND _06173_ _03108_ keymem.key_mem\[5\]\[56\] _06179_ sky130_fd_sc_hd__mux2_2
XFILLER_0_32_723 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_210_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_241_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24154_ VGND VPWR VPWR VGND clk _00647_ reset_n keymem.key_mem\[11\]\[19\] sky130_fd_sc_hd__dfrtp_2
X_21366_ VGND VPWR VPWR VGND _06140_ _02660_ keymem.key_mem\[5\]\[23\] _06143_ sky130_fd_sc_hd__mux2_2
XFILLER_0_32_778 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Right_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23105_ VGND VPWR VGND VPWR _07030_ _03449_ _06890_ _03451_ _07011_ sky130_fd_sc_hd__a211o_2
X_20317_ VGND VPWR _00928_ _05584_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24085_ VGND VPWR VPWR VGND clk _00578_ reset_n keymem.key_mem\[12\]\[78\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_31_299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21297_ VGND VPWR VPWR VGND _06098_ _03620_ keymem.key_mem\[6\]\[120\] _06105_ sky130_fd_sc_hd__mux2_2
X_23036_ VGND VPWR VGND VPWR _06987_ _03794_ _03215_ _06988_ sky130_fd_sc_hd__a21o_2
XFILLER_0_120_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_263_607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20248_ VGND VPWR _05548_ _10913_ _00895_ _05532_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_60_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20179_ VGND VPWR VPWR VGND _05504_ _03550_ keymem.key_mem\[10\]\[109\] _05510_ sky130_fd_sc_hd__mux2_2
X_24987_ VGND VPWR VPWR VGND clk _01480_ reset_n keymem.key_mem\[5\]\[84\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14740_ VPWR VGND VGND VPWR _09069_ _09103_ _09168_ _09138_ _10206_ _10205_ sky130_fd_sc_hd__o221a_2
XFILLER_0_58_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23938_ VGND VPWR VPWR VGND clk _00431_ reset_n keymem.key_mem\[13\]\[59\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_235_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11952_ VPWR VGND VGND VPWR _07554_ _07555_ _07530_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_42_Right_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14671_ VGND VPWR VGND VPWR _09368_ _10135_ _10137_ _10136_ _10138_ sky130_fd_sc_hd__o22a_2
X_11883_ VGND VPWR result[108] _07505_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23869_ VGND VPWR VPWR VGND clk _00362_ reset_n enc_block.block_w2_reg\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_1158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16410_ VGND VPWR VGND VPWR _02562_ _02571_ _02572_ _02556_ _02566_ sky130_fd_sc_hd__nor4_2
XFILLER_0_19_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13622_ VPWR VGND VPWR VGND _09031_ _09027_ _09017_ _08958_ _09094_ sky130_fd_sc_hd__or4_2
X_25608_ VGND VPWR VPWR VGND clk _02101_ reset_n keymem.key_mem\[0\]\[65\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_170_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17390_ VPWR VGND VGND VPWR _03476_ key[226] _09522_ sky130_fd_sc_hd__nand2_2
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16341_ VGND VPWR VGND VPWR _11250_ _11284_ _11464_ _11311_ _02504_ sky130_fd_sc_hd__o22a_2
XFILLER_0_27_517 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13553_ VGND VPWR VGND VPWR enc_block.block_w1_reg\[0\] _08948_ _09022_ _09023_ _09025_
+ _09024_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_54_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25539_ VGND VPWR VPWR VGND clk _02032_ reset_n keymem.key_mem\[1\]\[124\] sky130_fd_sc_hd__dfrtp_2
X_12504_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[35\] _07568_ keymem.key_mem\[6\]\[35\]
+ _07656_ _08072_ sky130_fd_sc_hd__a22o_2
XFILLER_0_183_179 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19060_ VGND VPWR VGND VPWR _04882_ keymem.key_mem_we _09725_ _04878_ _00373_ sky130_fd_sc_hd__a31o_2
X_16272_ VGND VPWR _11246_ _11412_ _02436_ _11278_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_13484_ VGND VPWR _08956_ _08955_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_129_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15223_ VGND VPWR VGND VPWR _10480_ _10475_ _10593_ _10508_ _10686_ sky130_fd_sc_hd__o22a_2
XFILLER_0_35_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_205_Left_472 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18011_ VGND VPWR VGND VPWR _03737_ keymem.prev_key1_reg\[127\] _03939_ _03738_ sky130_fd_sc_hd__a21oi_2
X_12435_ VGND VPWR _08009_ _07618_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_191_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_51_Right_51 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_129_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15154_ VGND VPWR _10618_ _10559_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_26_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12366_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[23\] _07582_ keymem.key_mem\[8\]\[23\]
+ _07539_ _07946_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_778 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_205_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14105_ VGND VPWR _09576_ _09431_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_240_1023 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_181_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15085_ VGND VPWR VGND VPWR _10510_ _10546_ _10519_ _10535_ _10549_ sky130_fd_sc_hd__o22a_2
X_19962_ VGND VPWR VPWR VGND _05389_ _10284_ keymem.key_mem\[10\]\[6\] _05396_ sky130_fd_sc_hd__mux2_2
X_12297_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[17\] _07645_ _07882_ _07875_ _07883_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_238_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18913_ VPWR VGND VPWR VGND _04752_ _04664_ _04751_ enc_block.block_w2_reg\[16\]
+ _04709_ _00356_ sky130_fd_sc_hd__a221o_2
X_14036_ VPWR VGND _09508_ _09507_ keymem.prev_key0_reg\[96\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_205_1198 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19893_ VGND VPWR VPWR VGND _05350_ keymem.key_mem\[11\]\[103\] _03511_ _05358_ sky130_fd_sc_hd__mux2_2
XFILLER_0_142_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_129_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18844_ VGND VPWR VGND VPWR _04689_ _04690_ _04600_ _04691_ enc_block.block_w2_reg\[9\]
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_235_832 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_214_Left_481 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_175_1220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18775_ VGND VPWR _04628_ enc_block.block_w1_reg\[7\] _04627_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_250_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_60_Right_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_89_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15987_ VGND VPWR _09512_ key[16] _11443_ _09987_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_37_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17726_ VPWR VGND VPWR VGND _02836_ _03750_ keymem.prev_key0_reg\[30\] _03730_ _00171_
+ sky130_fd_sc_hd__a22o_2
X_14938_ VGND VPWR _10402_ _08954_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_37_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_209_Right_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17657_ VGND VPWR VPWR VGND _03681_ _03700_ keymem.prev_key0_reg\[11\] _03701_ sky130_fd_sc_hd__mux2_2
X_14869_ VPWR VGND VGND VPWR _09641_ _09848_ _09825_ _10333_ _10334_ sky130_fd_sc_hd__and4b_2
X_16608_ VGND VPWR _02765_ _02764_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_147_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17588_ VGND VPWR VPWR VGND _03593_ keymem.key_mem\[14\]\[124\] _03647_ _03648_ sky130_fd_sc_hd__mux2_2
XFILLER_0_212_1158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_46_826 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19327_ VPWR VGND keymem.key_mem_we _05045_ _03533_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16539_ VGND VPWR VGND VPWR _11532_ keymem.rcon_logic.tmp_rcon\[2\] _02698_ _11502_
+ sky130_fd_sc_hd__nand3_2
XFILLER_0_70_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_223_Left_490 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19258_ VGND VPWR VGND VPWR _05001_ keymem.key_mem_we _03330_ _04999_ _00452_ sky130_fd_sc_hd__a31o_2
XFILLER_0_2_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_147_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18209_ VPWR VGND _04118_ enc_block.block_w2_reg\[12\] enc_block.block_w3_reg\[4\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_170_330 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_115_257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19189_ VPWR VGND keymem.key_mem\[13\]\[53\] _04960_ _04915_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_48_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21220_ VGND VPWR _01351_ _06064_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_218_Right_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_108_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_223_1221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_935 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_586 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21151_ VGND VPWR _01318_ _06028_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_160_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20102_ VGND VPWR VPWR VGND _05469_ _03259_ keymem.key_mem\[10\]\[72\] _05470_ sky130_fd_sc_hd__mux2_2
X_21082_ VGND VPWR _01285_ _05992_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20033_ VGND VPWR _00795_ _05433_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24910_ VGND VPWR VPWR VGND clk _01403_ reset_n keymem.key_mem\[5\]\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_186_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24841_ VGND VPWR VPWR VGND clk _01334_ reset_n keymem.key_mem\[6\]\[66\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_158_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_119_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_227_Right_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24772_ VGND VPWR VPWR VGND clk _01265_ reset_n keymem.key_mem\[7\]\[125\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_59_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21984_ VPWR VGND keymem.key_mem\[3\]\[56\] _06472_ _06469_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_119_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23723_ keymem.prev_key0_reg\[79\] clk _00220_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20935_ VGND VPWR VPWR VGND _05912_ _04995_ keymem.key_mem\[7\]\[77\] _05914_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_1_Right_797 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23654_ keymem.prev_key0_reg\[10\] clk _00151_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20866_ VGND VPWR VPWR VGND _05867_ _04945_ keymem.key_mem\[7\]\[45\] _05877_ sky130_fd_sc_hd__mux2_2
XFILLER_0_165_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22605_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[115\] _06777_ _06776_ _05064_ _02023_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_49_697 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23585_ VGND VPWR VPWR VGND clk _00086_ reset_n keymem.key_mem\[14\]\[74\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_165_157 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20797_ VPWR VGND keymem.key_mem\[7\]\[13\] _05840_ _05830_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_64_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25324_ VGND VPWR VPWR VGND clk _01817_ reset_n keymem.key_mem\[2\]\[37\] sky130_fd_sc_hd__dfrtp_2
X_22536_ VGND VPWR _06756_ _06701_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_228_1110 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_106_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25255_ VGND VPWR VPWR VGND clk _01748_ reset_n keymem.key_mem\[3\]\[96\] sky130_fd_sc_hd__dfrtp_2
X_22467_ VGND VPWR VPWR VGND _06726_ keymem.key_mem\[1\]\[27\] _02765_ _06728_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_594 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24206_ VGND VPWR VPWR VGND clk _00699_ reset_n keymem.key_mem\[11\]\[71\] sky130_fd_sc_hd__dfrtp_2
X_12220_ VGND VPWR _07811_ _07613_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21418_ VGND VPWR VPWR VGND _06162_ _03035_ keymem.key_mem\[5\]\[48\] _06170_ sky130_fd_sc_hd__mux2_2
XFILLER_0_66_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25186_ VGND VPWR VPWR VGND clk _01679_ reset_n keymem.key_mem\[3\]\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22398_ VGND VPWR _01903_ _06690_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_206_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12151_ VGND VPWR VGND VPWR _07747_ _07743_ keymem.key_mem\[10\]\[7\] _07745_ _07746_
+ sky130_fd_sc_hd__a211o_2
X_24137_ VGND VPWR VPWR VGND clk _00630_ reset_n keymem.key_mem\[11\]\[2\] sky130_fd_sc_hd__dfrtp_2
X_21349_ VGND VPWR VPWR VGND _06128_ _11148_ keymem.key_mem\[5\]\[15\] _06134_ sky130_fd_sc_hd__mux2_2
XFILLER_0_27_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24068_ VGND VPWR VPWR VGND clk _00561_ reset_n keymem.key_mem\[12\]\[61\] sky130_fd_sc_hd__dfrtp_2
X_12082_ VPWR VGND VPWR VGND _07680_ keymem.key_mem\[3\]\[4\] _07602_ keymem.key_mem\[10\]\[4\]
+ _07560_ _07681_ sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_71_1_Left_338 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15910_ _11340_ _11366_ _11222_ _11365_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_23019_ VGND VPWR VPWR VGND _06960_ _06978_ keymem.prev_key1_reg\[59\] _06979_ sky130_fd_sc_hd__mux2_2
X_16890_ VGND VPWR _00059_ _03026_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15841_ VGND VPWR VPWR VGND _11173_ _11247_ _11233_ _11297_ sky130_fd_sc_hd__or3_2
XFILLER_0_95_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_164_2_Left_635 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_137_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18560_ VGND VPWR _04435_ enc_block.block_w3_reg\[12\] enc_block.block_w0_reg\[4\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15772_ VGND VPWR _11228_ _11197_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12984_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[82\] _07818_ keymem.key_mem\[9\]\[82\]
+ _07705_ _08505_ sky130_fd_sc_hd__a22o_2
X_17511_ VGND VPWR VPWR VGND _03534_ keymem.key_mem\[14\]\[114\] _03580_ _03581_ sky130_fd_sc_hd__mux2_2
XFILLER_0_8_1029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11935_ VPWR VGND VGND VPWR _07537_ _07538_ _07527_ sky130_fd_sc_hd__nor2_2
X_14723_ VPWR VGND VGND VPWR _10190_ keylen _09927_ sky130_fd_sc_hd__nand2_2
X_18491_ VPWR VGND _04373_ enc_block.block_w0_reg\[5\] enc_block.block_w1_reg\[29\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_217_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14654_ VPWR VGND VGND VPWR _09311_ _09378_ _10121_ _09443_ _09396_ sky130_fd_sc_hd__o22ai_2
X_17442_ VGND VPWR VGND VPWR _03521_ _10328_ _02877_ key[105] sky130_fd_sc_hd__o21a_2
X_11866_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[4\] dec_new_block\[100\]
+ _07497_ sky130_fd_sc_hd__mux2_2
XFILLER_0_262_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_28_826 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13605_ VGND VPWR _09077_ _09076_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14585_ VPWR VGND VPWR VGND _09581_ _09784_ _10053_ _10052_ _09580_ sky130_fd_sc_hd__or4b_2
XFILLER_0_71_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17373_ VGND VPWR _00107_ _03461_ VPWR VGND sky130_fd_sc_hd__buf_1
X_11797_ VGND VPWR result[65] _07462_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_32_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19112_ VGND VPWR VGND VPWR _04911_ keymem.key_mem_we _02689_ _04908_ _00396_ sky130_fd_sc_hd__a31o_2
XFILLER_0_171_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_144_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_347 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13536_ VGND VPWR VGND VPWR _09008_ _08953_ _08950_ keymem.prev_key1_reg\[2\] _08969_
+ _08964_ sky130_fd_sc_hd__a32o_2
X_16324_ VGND VPWR VPWR VGND _10993_ _11018_ _02485_ _02487_ sky130_fd_sc_hd__or3_2
XFILLER_0_137_371 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16255_ VGND VPWR _11323_ _11236_ _02419_ _11473_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_19043_ VGND VPWR _04868_ enc_block.block_w3_reg\[23\] enc_block.block_w1_reg\[7\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_881 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13467_ VPWR VGND VPWR VGND enc_block.sword_ctr_inc _08939_ enc_block.enc_ctrl_reg\[3\]
+ enc_block.enc_ctrl_reg\[2\] sky130_fd_sc_hd__or3b_2
X_15206_ VGND VPWR VGND VPWR _10667_ _10538_ _10528_ _10668_ _10669_ sky130_fd_sc_hd__o22a_2
XFILLER_0_242_1107 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12418_ VGND VPWR enc_block.round_key\[27\] _07993_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_211_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16186_ VPWR VGND VGND VPWR _11473_ _02351_ _11219_ sky130_fd_sc_hd__nor2_2
XFILLER_0_23_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13398_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[123\] _07583_ keymem.key_mem\[9\]\[123\]
+ _07592_ _08878_ sky130_fd_sc_hd__a22o_2
XFILLER_0_112_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15137_ VPWR VGND VPWR VGND _10483_ _10409_ _10452_ _10412_ _10601_ sky130_fd_sc_hd__or4_2
XFILLER_0_11_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12349_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[21\] _07608_ keymem.key_mem\[14\]\[21\]
+ _07582_ _07931_ sky130_fd_sc_hd__a22o_2
XFILLER_0_199_1039 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_142_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15068_ VPWR VGND VPWR VGND _10525_ _10531_ _10532_ _10517_ _10523_ sky130_fd_sc_hd__or4b_2
X_19945_ _07387_ _05385_ keymem.key_mem_we keymem.round_ctr_reg\[1\] VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__and3_2
XFILLER_0_103_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_120_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_821 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14019_ VGND VPWR VGND VPWR _09341_ _09302_ _09336_ _09419_ _09491_ sky130_fd_sc_hd__o22a_2
XFILLER_0_177_1315 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19876_ VGND VPWR VPWR VGND _05339_ keymem.key_mem\[11\]\[95\] _03460_ _05349_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_96_2_Left_567 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_177_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18827_ VGND VPWR _04675_ enc_block.block_w0_reg\[15\] _04592_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_120_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_235_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18758_ VGND VPWR _04613_ _04599_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17709_ VGND VPWR VGND VPWR _03737_ keymem.prev_key1_reg\[25\] _03739_ _03738_ sky130_fd_sc_hd__a21oi_2
X_18689_ VPWR VGND VGND VPWR _04512_ _04551_ _04256_ sky130_fd_sc_hd__nor2_2
XFILLER_0_77_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20720_ VGND VPWR _01119_ _05796_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_187_260 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_37_1186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20651_ VPWR VGND VGND VPWR _05676_ _05760_ keymem.key_mem\[8\]\[75\] sky130_fd_sc_hd__nor2_2
XFILLER_0_92_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23370_ VGND VPWR VGND VPWR _07244_ _04266_ _07095_ _07245_ enc_block.block_w3_reg\[16\]
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_50_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20582_ VGND VPWR VPWR VGND _05714_ _02972_ keymem.key_mem\[8\]\[42\] _05724_ sky130_fd_sc_hd__mux2_2
XFILLER_0_188_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_103 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22321_ VGND VPWR _01866_ _06650_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_60_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_263 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_264_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25040_ VGND VPWR VPWR VGND clk _01533_ reset_n keymem.key_mem\[4\]\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_121_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22252_ VGND VPWR _01833_ _06614_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_564 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_60_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21203_ VPWR VGND VGND VPWR _06056_ keymem.key_mem\[6\]\[75\] _05985_ sky130_fd_sc_hd__nand2_2
X_22183_ VGND VPWR _06578_ _06553_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_2_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21134_ VGND VPWR VPWR VGND _06018_ _02972_ keymem.key_mem\[6\]\[42\] _06020_ sky130_fd_sc_hd__mux2_2
XFILLER_0_160_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21065_ VGND VPWR _05983_ _05971_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_258_1158 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_219_1109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_22_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20016_ VGND VPWR VPWR VGND _05424_ _02862_ keymem.key_mem\[10\]\[31\] _05425_ sky130_fd_sc_hd__mux2_2
XFILLER_0_195_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24824_ VGND VPWR VPWR VGND clk _01317_ reset_n keymem.key_mem\[6\]\[49\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_193_1161 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_225_194 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_154_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24755_ VGND VPWR VPWR VGND clk _01248_ reset_n keymem.key_mem\[7\]\[108\] sky130_fd_sc_hd__dfrtp_2
X_21967_ VGND VPWR VPWR VGND _06462_ _04950_ keymem.key_mem\[3\]\[48\] _06463_ sky130_fd_sc_hd__mux2_2
XFILLER_0_154_1167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_213_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11720_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[27\] dec_new_block\[27\]
+ _07424_ sky130_fd_sc_hd__mux2_2
X_23706_ keymem.prev_key0_reg\[62\] clk _00203_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20918_ VPWR VGND keymem.key_mem\[7\]\[69\] _05905_ _05899_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_189_1208 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24686_ VGND VPWR VPWR VGND clk _01179_ reset_n keymem.key_mem\[7\]\[39\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_132_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21898_ VGND VPWR VGND VPWR _06425_ keymem.key_mem_we _11447_ _06420_ _01668_ sky130_fd_sc_hd__a31o_2
XPHY_EDGE_ROW_180_2_Right_252 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23637_ VGND VPWR VPWR VGND clk _00138_ reset_n keymem.key_mem\[14\]\[126\] sky130_fd_sc_hd__dfrtp_2
X_11651_ VGND VPWR _07388_ keymem.round_ctr_reg\[2\] keylen VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20849_ VGND VPWR _01176_ _05868_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_132_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14370_ VPWR VGND VGND VPWR _09056_ _09019_ _09840_ _09132_ _09053_ sky130_fd_sc_hd__o22ai_2
X_23568_ VGND VPWR VPWR VGND clk _00069_ reset_n keymem.key_mem\[14\]\[57\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_382 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_119_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13321_ VPWR VGND VPWR VGND keymem.key_mem\[8\]\[115\] _07752_ keymem.key_mem\[1\]\[115\]
+ _07670_ _08809_ sky130_fd_sc_hd__a22o_2
X_25307_ VGND VPWR VPWR VGND clk _01800_ reset_n keymem.key_mem\[2\]\[20\] sky130_fd_sc_hd__dfrtp_2
X_22519_ VGND VPWR VPWR VGND _06739_ keymem.key_mem\[1\]\[60\] _03150_ _06747_ sky130_fd_sc_hd__mux2_2
X_23499_ VPWR VGND VPWR VGND _07359_ _07167_ _07357_ sky130_fd_sc_hd__or2_2
XFILLER_0_51_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16040_ VGND VPWR VGND VPWR _11236_ _11379_ _11473_ _11314_ _11495_ sky130_fd_sc_hd__o22a_2
X_25238_ VGND VPWR VPWR VGND clk _01731_ reset_n keymem.key_mem\[3\]\[79\] sky130_fd_sc_hd__dfrtp_2
X_13252_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[108\] _07984_ keymem.key_mem\[2\]\[108\]
+ _08131_ _08747_ sky130_fd_sc_hd__a22o_2
XFILLER_0_51_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_243_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_161_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12203_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[11\] _07568_ keymem.key_mem\[9\]\[11\]
+ _07592_ _07795_ sky130_fd_sc_hd__a22o_2
X_13183_ VGND VPWR VGND VPWR _08685_ _07839_ keymem.key_mem\[11\]\[101\] _08682_ _08684_
+ sky130_fd_sc_hd__a211o_2
X_25169_ VGND VPWR VPWR VGND clk _01662_ reset_n keymem.key_mem\[3\]\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_62_1246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12134_ VGND VPWR _07730_ _07667_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_209_607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_143_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17991_ VGND VPWR VGND VPWR _03926_ _03925_ _03675_ _03618_ sky130_fd_sc_hd__and3b_2
XFILLER_0_40_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19730_ VGND VPWR VPWR VGND _05270_ keymem.key_mem\[11\]\[25\] _02721_ _05273_ sky130_fd_sc_hd__mux2_2
X_16942_ VGND VPWR VPWR VGND _03072_ _02475_ _03074_ _02496_ _03073_ sky130_fd_sc_hd__o211a_2
X_12065_ VGND VPWR _07665_ _07552_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_19_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_779 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19661_ VGND VPWR _00622_ _05234_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16873_ VGND VPWR VPWR VGND _09521_ key[174] keymem.prev_key1_reg\[46\] _03011_ sky130_fd_sc_hd__mux2_2
XFILLER_0_216_150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18612_ VGND VPWR _04482_ _04480_ _04481_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15824_ VGND VPWR _11280_ _11279_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19592_ VGND VPWR _00589_ _05198_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_232_654 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_220_805 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18543_ VGND VPWR VGND VPWR _04419_ _04418_ _04420_ _03966_ sky130_fd_sc_hd__a21oi_2
X_15755_ VGND VPWR _11211_ _11210_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12967_ VGND VPWR VGND VPWR _07984_ keymem.key_mem\[14\]\[80\] _08487_ _08489_ _08490_
+ _07662_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_231_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_172_1278 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11918_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[30\] dec_new_block\[126\]
+ _07523_ sky130_fd_sc_hd__mux2_2
X_14706_ VPWR VGND VGND VPWR _09110_ _10173_ _09174_ sky130_fd_sc_hd__nor2_2
XFILLER_0_129_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_206_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18474_ VPWR VGND VGND VPWR _04358_ _04353_ _04356_ sky130_fd_sc_hd__nand2_2
XFILLER_0_47_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15686_ VGND VPWR VPWR VGND keymem.round_ctr_reg\[0\] _11142_ _11104_ _11143_ sky130_fd_sc_hd__mux2_2
XFILLER_0_129_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12898_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[73\] _07730_ keymem.key_mem\[9\]\[73\]
+ _07705_ _08428_ sky130_fd_sc_hd__a22o_2
XFILLER_0_142_14 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_74_206 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_150_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17425_ VGND VPWR VPWR VGND _03467_ keymem.key_mem\[14\]\[102\] _03506_ _03507_ sky130_fd_sc_hd__mux2_2
X_11849_ VGND VPWR result[91] _07488_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14637_ VPWR VGND VGND VPWR _09353_ _10104_ _09341_ sky130_fd_sc_hd__nor2_2
XFILLER_0_111_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_200_573 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_142_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_7_517 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_248_1327 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14568_ VGND VPWR VGND VPWR _09392_ _09487_ _09420_ _09475_ _10036_ sky130_fd_sc_hd__o22a_2
XFILLER_0_129_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17356_ VPWR VGND VPWR VGND _03446_ keymem.prev_key0_reg\[94\] sky130_fd_sc_hd__inv_2
X_16307_ VGND VPWR VGND VPWR _10960_ _10948_ keymem.prev_key1_reg\[116\] _02471_ sky130_fd_sc_hd__a21o_2
XFILLER_0_3_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13519_ VGND VPWR _08991_ _08990_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14499_ VGND VPWR VGND VPWR _09107_ _09154_ _09122_ _09160_ _09968_ sky130_fd_sc_hd__o22a_2
X_17287_ VGND VPWR VPWR VGND _03384_ keymem.key_mem\[14\]\[86\] _03383_ _03385_ sky130_fd_sc_hd__mux2_2
XFILLER_0_261_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19026_ VPWR VGND VPWR VGND _04853_ _04788_ _04852_ enc_block.block_w2_reg\[28\]
+ _04613_ _00368_ sky130_fd_sc_hd__a221o_2
XFILLER_0_109_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16238_ VGND VPWR _02403_ keymem.prev_key1_reg\[83\] _02402_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_261_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16169_ VPWR VGND VPWR VGND _11622_ _11623_ _09932_ _11561_ sky130_fd_sc_hd__or3b_2
XFILLER_0_224_1393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_259_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19928_ VGND VPWR _00747_ _05376_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_43_1190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_255_Right_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19859_ VGND VPWR _00714_ _05340_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_235_470 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_183_10 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_78_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22870_ VGND VPWR VGND VPWR _02179_ _06886_ _06882_ keymem.prev_key1_reg\[2\] sky130_fd_sc_hd__o21a_2
XFILLER_0_190_1323 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_190_1345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21821_ VGND VPWR _01634_ _06382_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_890 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24540_ VGND VPWR VPWR VGND clk _01033_ reset_n keymem.key_mem\[8\]\[21\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_190_1389 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21752_ VGND VPWR _01601_ _06346_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_231_1353 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20703_ VGND VPWR _01111_ _05787_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24471_ VGND VPWR VPWR VGND clk _00964_ reset_n keymem.key_mem\[9\]\[80\] sky130_fd_sc_hd__dfrtp_2
X_21683_ VGND VPWR _01568_ _06310_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_58_280 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23422_ VPWR VGND _07291_ _07140_ enc_block.block_w3_reg\[30\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_114_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20634_ VGND VPWR _01078_ _05751_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_11_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23353_ VGND VPWR VPWR VGND _07093_ enc_block.block_w3_reg\[14\] _04135_ _07230_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_6_550 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20565_ VGND VPWR _01045_ _05715_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_184_1149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_6_583 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22304_ VGND VPWR _01858_ _06641_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_190_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23284_ VGND VPWR _07167_ enc_block.block_w2_reg\[7\] enc_block.block_w1_reg\[15\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_166_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_85_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20496_ VGND VPWR _01013_ _05678_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_264_1195 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_260_1037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25023_ VGND VPWR VPWR VGND clk _01516_ reset_n keymem.key_mem\[5\]\[120\] sky130_fd_sc_hd__dfrtp_2
X_22235_ VGND VPWR _01825_ _06605_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_383 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22166_ VGND VPWR _01792_ _06569_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_125_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_160_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21117_ VGND VPWR VPWR VGND _06007_ _02893_ keymem.key_mem\[6\]\[34\] _06011_ sky130_fd_sc_hd__mux2_2
XFILLER_0_22_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22097_ VGND VPWR _01761_ _06531_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_96_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_121_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21048_ VGND VPWR _01269_ _05974_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_156_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_100_1_Right_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_227_993 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_254_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13870_ VGND VPWR VPWR VGND _09261_ _09315_ _09254_ _09342_ sky130_fd_sc_hd__or3_2
XFILLER_0_96_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_236_1253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_92_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12821_ VGND VPWR enc_block.round_key\[65\] _08358_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24807_ VGND VPWR VPWR VGND clk _01300_ reset_n keymem.key_mem\[6\]\[32\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_201_304 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_838 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22999_ VGND VPWR VPWR VGND _06960_ _06966_ keymem.prev_key1_reg\[51\] _06967_ sky130_fd_sc_hd__mux2_2
X_25787_ keymem.prev_key1_reg\[103\] clk _02280_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_9_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15540_ VPWR VGND VPWR VGND _10996_ _10998_ _10997_ _10919_ _10999_ sky130_fd_sc_hd__or4_2
X_12752_ VGND VPWR enc_block.round_key\[58\] _08296_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_243_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24738_ VGND VPWR VPWR VGND clk _01231_ reset_n keymem.key_mem\[7\]\[91\] sky130_fd_sc_hd__dfrtp_2
X_11703_ VGND VPWR result[18] _07415_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_210_1415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15471_ VPWR VGND VGND VPWR _10536_ _10931_ _10565_ sky130_fd_sc_hd__nor2_2
XFILLER_0_132_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12683_ VGND VPWR VGND VPWR _07841_ keymem.key_mem\[4\]\[52\] _08231_ _08233_ _08234_
+ _08069_ sky130_fd_sc_hd__a2111o_2
X_24669_ VGND VPWR VPWR VGND clk _01162_ reset_n keymem.key_mem\[7\]\[22\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_181_2_Right_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14422_ VGND VPWR VGND VPWR _09891_ _09444_ _09358_ _09487_ _09392_ _09890_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_132_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17210_ VGND VPWR _00090_ _03315_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_33_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11634_ VGND VPWR _07374_ _07373_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_167_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18190_ VPWR VGND VGND VPWR _04100_ _04101_ _04098_ sky130_fd_sc_hd__nor2_2
XFILLER_0_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14353_ VPWR VGND VGND VPWR _09113_ _09121_ _09823_ _09173_ _09148_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_64_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17141_ VGND VPWR _00083_ _03253_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_167_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13304_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[113\] _08714_ _08793_ _08789_ _08794_
+ sky130_fd_sc_hd__o22a_2
X_17072_ VGND VPWR VGND VPWR _03189_ _03191_ _03188_ keylen _03192_ sky130_fd_sc_hd__a2bb2o_2
X_14284_ VPWR VGND VGND VPWR _09754_ _09303_ _09304_ sky130_fd_sc_hd__nand2_2
XFILLER_0_12_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16023_ _11477_ _11478_ _11224_ _11290_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_122_355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_243_1257 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13235_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[106\] _08714_ _08731_ _08727_ _08732_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_27_1130 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13166_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[100\] _07629_ keymem.key_mem\[12\]\[100\]
+ _07579_ _08669_ sky130_fd_sc_hd__a22o_2
XFILLER_0_104_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_375 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_62_1087 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_196_1009 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_143_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12117_ VGND VPWR _07714_ _07556_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_104_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17974_ VGND VPWR _00255_ _03914_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13097_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[93\] _07872_ keymem.key_mem\[6\]\[93\]
+ _07639_ _08607_ sky130_fd_sc_hd__a22o_2
XFILLER_0_40_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19713_ VGND VPWR VPWR VGND _05259_ keymem.key_mem\[11\]\[17\] _11547_ _05264_ sky130_fd_sc_hd__mux2_2
XFILLER_0_100_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16925_ VPWR VGND VPWR VGND _02396_ _03058_ _09932_ _02399_ sky130_fd_sc_hd__or3b_2
X_12048_ VGND VPWR _07648_ _07647_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_40_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1028 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_178_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19644_ VGND VPWR _00614_ _05225_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16856_ VPWR VGND VPWR VGND keylen _02995_ _02994_ _10968_ _02993_ _02996_ sky130_fd_sc_hd__a221o_2
XFILLER_0_232_440 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_75_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15807_ VGND VPWR _11263_ _11233_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19575_ VGND VPWR VPWR VGND _05183_ _05002_ keymem.key_mem\[12\]\[81\] _05190_ sky130_fd_sc_hd__mux2_2
X_16787_ VGND VPWR VPWR VGND _10277_ _02930_ _02933_ _02496_ _02932_ sky130_fd_sc_hd__o211a_2
X_13999_ VGND VPWR VPWR VGND _09462_ _09470_ _09457_ _09471_ sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_159_1_Left_426 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18526_ VPWR VGND VPWR VGND _04404_ block[73] _04330_ enc_block.block_w3_reg\[9\]
+ _04276_ _04405_ sky130_fd_sc_hd__a221o_2
XFILLER_0_246_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15738_ VGND VPWR VGND VPWR _11194_ enc_block.block_w2_reg\[20\] enc_block.sword_ctr_reg\[1\]
+ enc_block.sword_ctr_reg\[0\] sky130_fd_sc_hd__and3b_2
XFILLER_0_220_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1061 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_150_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18457_ VPWR VGND _04342_ enc_block.block_w1_reg\[27\] enc_block.block_w2_reg\[19\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_115_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15669_ VGND VPWR VPWR VGND _11126_ _10953_ _10619_ _10572_ _10714_ sky130_fd_sc_hd__o31a_2
XFILLER_0_111_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17408_ VGND VPWR VGND VPWR _03491_ _03488_ _03492_ _03490_ sky130_fd_sc_hd__nand3_2
XFILLER_0_150_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18388_ VPWR VGND VPWR VGND _04280_ block[125] _04213_ enc_block.block_w0_reg\[29\]
+ _04276_ _04281_ sky130_fd_sc_hd__a221o_2
XFILLER_0_189_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_347 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_55_250 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_111_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17339_ VGND VPWR VGND VPWR key[92] _09930_ _03430_ _03429_ _03431_ sky130_fd_sc_hd__o22a_2
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_86_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20350_ VGND VPWR _00944_ _05601_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_15_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_629 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19009_ VPWR VGND _04838_ enc_block.block_w1_reg\[3\] enc_block.block_w3_reg\[18\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_261_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_140_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20281_ VGND VPWR _00911_ _05565_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_11_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_113_388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22020_ VPWR VGND keymem.key_mem\[3\]\[73\] _06491_ _06484_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_144_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23971_ VGND VPWR VPWR VGND clk _00464_ reset_n keymem.key_mem\[13\]\[92\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_1565 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_157_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_192_1418 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_93_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22922_ VGND VPWR VGND VPWR _02596_ _06890_ _02606_ _06919_ sky130_fd_sc_hd__a21o_2
X_25710_ keymem.prev_key1_reg\[26\] clk _02203_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_93_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_602 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25641_ VGND VPWR VPWR VGND clk _02134_ reset_n keymem.key_mem\[0\]\[98\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_211_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22853_ VGND VPWR VGND VPWR _06875_ _06874_ _05818_ keymem.round_ctr_rst sky130_fd_sc_hd__and3b_2
XFILLER_0_233_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_196_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_52_1201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21804_ VGND VPWR _01626_ _06373_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25572_ VGND VPWR VPWR VGND clk _02065_ reset_n keymem.key_mem\[0\]\[29\] sky130_fd_sc_hd__dfrtp_2
X_22784_ VGND VPWR VPWR VGND _06784_ keymem.key_mem\[0\]\[91\] _03427_ _06853_ sky130_fd_sc_hd__mux2_2
XFILLER_0_211_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24523_ VGND VPWR VPWR VGND clk _01016_ reset_n keymem.key_mem\[8\]\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_133_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21735_ VGND VPWR _01593_ _06337_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_231_1172 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24454_ VGND VPWR VPWR VGND clk _00947_ reset_n keymem.key_mem\[9\]\[63\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_80_1_Left_347 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21666_ VGND VPWR _01560_ _06301_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23405_ VGND VPWR _07276_ enc_block.block_w2_reg\[4\] enc_block.block_w1_reg\[12\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_163_244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20617_ VGND VPWR _01070_ _05742_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24385_ VGND VPWR VPWR VGND clk _00878_ reset_n keymem.key_mem\[10\]\[122\] sky130_fd_sc_hd__dfrtp_2
X_21597_ VGND VPWR _01527_ _06265_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23336_ VPWR VGND VPWR VGND _07214_ enc_block.block_w2_reg\[4\] enc_block.block_w2_reg\[5\]
+ sky130_fd_sc_hd__or2_2
XFILLER_0_244_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20548_ VGND VPWR _01037_ _05706_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_173_2_Left_644 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_692 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23267_ VPWR VGND VGND VPWR _07152_ _07148_ _07150_ sky130_fd_sc_hd__nand2_2
XFILLER_0_244_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20479_ VGND VPWR VPWR VGND _05660_ _03633_ keymem.key_mem\[9\]\[122\] _05669_ sky130_fd_sc_hd__mux2_2
X_13020_ VPWR VGND VPWR VGND _08537_ keymem.key_mem\[11\]\[85\] _08090_ keymem.key_mem\[2\]\[85\]
+ _07733_ _08538_ sky130_fd_sc_hd__a221o_2
X_25006_ VGND VPWR VPWR VGND clk _01499_ reset_n keymem.key_mem\[5\]\[103\] sky130_fd_sc_hd__dfrtp_2
X_22218_ VGND VPWR _01817_ _06596_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23198_ VPWR VGND VGND VPWR _07088_ _07089_ _03966_ sky130_fd_sc_hd__nor2_2
XFILLER_0_140_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22149_ VGND VPWR VPWR VGND _06554_ _10193_ keymem.key_mem\[2\]\[5\] _06560_ sky130_fd_sc_hd__mux2_2
XFILLER_0_101_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1285 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_140_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14971_ VGND VPWR VGND VPWR _10435_ _10434_ _10433_ keymem.prev_key1_reg\[15\] _09003_
+ _09002_ sky130_fd_sc_hd__a32o_2
XFILLER_0_101_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_238_1348 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_22_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16710_ VGND VPWR VPWR VGND _02662_ keymem.key_mem\[14\]\[31\] _02862_ _02863_ sky130_fd_sc_hd__mux2_2
X_13922_ VPWR VGND VPWR VGND _09385_ _09393_ _09394_ _09359_ _09369_ sky130_fd_sc_hd__or4b_2
X_17690_ VGND VPWR _03723_ _03674_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_1_Right_702 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_96_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16641_ VGND VPWR _02796_ _02793_ _02795_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_13853_ VPWR VGND VPWR VGND _09325_ _09313_ _09324_ sky130_fd_sc_hd__or2_2
X_25839_ VGND VPWR VPWR VGND clk _02332_ reset_n enc_block.block_w3_reg\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_251_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12804_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[64\] _08032_ keymem.key_mem\[12\]\[64\]
+ _07621_ _08343_ sky130_fd_sc_hd__a22o_2
X_19360_ VGND VPWR VPWR VGND _05067_ _05066_ keymem.key_mem\[13\]\[116\] _05068_ sky130_fd_sc_hd__mux2_2
X_16572_ VGND VPWR _02730_ keymem.prev_key0_reg\[26\] _02729_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_13784_ enc_block.sword_ctr_reg\[1\] _09256_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[26\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_18311_ VPWR VGND VGND VPWR _04211_ _04212_ _04190_ sky130_fd_sc_hd__nor2_2
X_15523_ VGND VPWR VGND VPWR _10535_ _10574_ _10646_ _10462_ _10981_ _10982_ sky130_fd_sc_hd__o32a_2
X_19291_ VPWR VGND keymem.key_mem_we _05021_ _03452_ VPWR VGND sky130_fd_sc_hd__and2_2
X_12735_ VPWR VGND VPWR VGND _08280_ keymem.key_mem\[13\]\[57\] _07835_ keymem.key_mem\[8\]\[57\]
+ _07753_ _08281_ sky130_fd_sc_hd__a221o_2
X_18242_ VGND VPWR _04149_ _04148_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_44_209 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12666_ VPWR VGND VPWR VGND _08218_ keymem.key_mem\[14\]\[50\] _07706_ keymem.key_mem\[2\]\[50\]
+ _07733_ _08219_ sky130_fd_sc_hd__a221o_2
X_15454_ VGND VPWR _10914_ _09541_ _00023_ _10913_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_182_2_Right_254 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14405_ VGND VPWR VGND VPWR _09312_ _09450_ _09576_ _09873_ _09874_ sky130_fd_sc_hd__o22a_2
X_18173_ VPWR VGND VGND VPWR _04086_ _04004_ _04085_ sky130_fd_sc_hd__nand2_2
X_15385_ VGND VPWR _10845_ _10667_ _10846_ _10455_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_12597_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[44\] _07969_ keymem.key_mem\[2\]\[44\]
+ _07733_ _08156_ sky130_fd_sc_hd__a22o_2
XFILLER_0_0_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_68_1252 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_119 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17124_ _10263_ _03238_ _03237_ _10264_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_14336_ VPWR VGND VPWR VGND _09806_ _09113_ _09082_ sky130_fd_sc_hd__or2_2
XFILLER_0_29_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_107_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1199 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14267_ VGND VPWR VGND VPWR _09737_ _09443_ _09403_ _09311_ sky130_fd_sc_hd__o21a_2
XFILLER_0_52_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_122_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17055_ VPWR VGND VPWR VGND _03176_ key[63] _09719_ sky130_fd_sc_hd__or2_2
XFILLER_0_0_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_110_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16006_ VGND VPWR VGND VPWR _11236_ _11336_ _11460_ _11404_ _11461_ sky130_fd_sc_hd__o22a_2
X_13218_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[105\] _07656_ keymem.key_mem\[11\]\[105\]
+ _07658_ _08716_ sky130_fd_sc_hd__a22o_2
XFILLER_0_0_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14198_ VPWR VGND VPWR VGND _09664_ _09668_ _09669_ _09662_ _09663_ sky130_fd_sc_hd__or4b_2
XFILLER_0_237_521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_695 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13149_ VGND VPWR VGND VPWR _07842_ keymem.key_mem\[9\]\[98\] _08651_ _08653_ _08654_
+ _08599_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_196_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_554 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_104_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17957_ VGND VPWR VPWR VGND _03896_ _03902_ keymem.prev_key0_reg\[109\] _03903_ sky130_fd_sc_hd__mux2_2
XFILLER_0_224_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16908_ VGND VPWR VPWR VGND _09511_ key[177] keymem.prev_key1_reg\[49\] _03043_ sky130_fd_sc_hd__mux2_2
XFILLER_0_224_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_75_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17888_ VGND VPWR VPWR VGND _03836_ _03855_ keymem.prev_key0_reg\[87\] _03856_ sky130_fd_sc_hd__mux2_2
XFILLER_0_139_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19627_ VGND VPWR VPWR VGND _05216_ _05045_ keymem.key_mem\[12\]\[106\] _05217_ sky130_fd_sc_hd__mux2_2
XFILLER_0_164_56 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16839_ VGND VPWR _10378_ keymem.prev_key1_reg\[43\] _02980_ keymem.prev_key1_reg\[75\]
+ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_221_922 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_75_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1183 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_220_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19558_ VGND VPWR VGND VPWR _05180_ keymem.key_mem_we _03268_ _05164_ _00573_ sky130_fd_sc_hd__a31o_2
XFILLER_0_250_1047 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_215_1189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18509_ VGND VPWR VGND VPWR _04388_ enc_block.round_key\[71\] _04149_ _04390_ sky130_fd_sc_hd__a21o_2
X_19489_ VGND VPWR VPWR VGND _05138_ _04937_ keymem.key_mem\[12\]\[41\] _05144_ sky130_fd_sc_hd__mux2_2
X_21520_ VGND VPWR _01492_ _06223_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_8_634 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_180_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_773 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_1216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_145_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21451_ VGND VPWR _01459_ _06187_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_44_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_266 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_12_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1255 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_43_242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20402_ VGND VPWR VPWR VGND _05627_ _03374_ keymem.key_mem\[9\]\[85\] _05629_ sky130_fd_sc_hd__mux2_2
XFILLER_0_86_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24170_ VGND VPWR VPWR VGND clk _00663_ reset_n keymem.key_mem\[11\]\[35\] sky130_fd_sc_hd__dfrtp_2
X_21382_ VGND VPWR _06151_ _06116_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_146_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_275 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_261_1121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_226_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23121_ VGND VPWR VPWR VGND _07032_ _07039_ keymem.prev_key1_reg\[100\] _07040_ sky130_fd_sc_hd__mux2_2
X_20333_ VGND VPWR VPWR VGND _05591_ _03075_ keymem.key_mem\[9\]\[52\] _05593_ sky130_fd_sc_hd__mux2_2
XFILLER_0_47_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1187 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23052_ VGND VPWR VGND VPWR _06888_ keymem.prev_key1_reg\[72\] _06998_ _02249_ sky130_fd_sc_hd__o21ba_2
X_20264_ VGND VPWR _00903_ _05556_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22003_ VGND VPWR VPWR VGND _06462_ _04975_ keymem.key_mem\[3\]\[65\] _06482_ sky130_fd_sc_hd__mux2_2
X_20195_ VGND VPWR _00872_ _05518_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_122_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_157_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_215_259 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23954_ VGND VPWR VPWR VGND clk _00447_ reset_n keymem.key_mem\[13\]\[75\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_760 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_157_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22905_ VGND VPWR VGND VPWR _02192_ _06908_ _06882_ keymem.prev_key1_reg\[15\] sky130_fd_sc_hd__o21a_2
XFILLER_0_212_933 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23885_ VGND VPWR VPWR VGND clk _00378_ reset_n keymem.key_mem\[13\]\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_19_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25624_ VGND VPWR VPWR VGND clk _02117_ reset_n keymem.key_mem\[0\]\[81\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_211_443 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22836_ VPWR VGND VGND VPWR _06861_ _06867_ _08922_ sky130_fd_sc_hd__nor2_2
XFILLER_0_6_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_334 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22767_ VGND VPWR _02116_ _06846_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_211_498 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25555_ VGND VPWR VPWR VGND clk _02048_ reset_n keymem.key_mem\[0\]\[12\] sky130_fd_sc_hd__dfrtp_2
X_12520_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[37\] _07845_ keymem.key_mem\[13\]\[37\]
+ _07834_ _08086_ sky130_fd_sc_hd__a22o_2
X_21718_ VGND VPWR _01585_ _06328_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24506_ VGND VPWR VPWR VGND clk _00999_ reset_n keymem.key_mem\[9\]\[115\] sky130_fd_sc_hd__dfrtp_2
X_25486_ VGND VPWR VPWR VGND clk _01979_ reset_n keymem.key_mem\[1\]\[71\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_136_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22698_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[39\] _06790_ _06789_ _04933_ _02075_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_47_570 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_168_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12451_ VPWR VGND VPWR VGND _08023_ keymem.key_mem\[14\]\[30\] _07706_ keymem.key_mem\[2\]\[30\]
+ _07733_ _08024_ sky130_fd_sc_hd__a221o_2
X_24437_ VGND VPWR VPWR VGND clk _00930_ reset_n keymem.key_mem\[9\]\[46\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_227_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21649_ VGND VPWR _01552_ _06292_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_30_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15170_ VPWR VGND VPWR VGND _10397_ _10466_ _10403_ _10392_ _10634_ sky130_fd_sc_hd__or4_2
XFILLER_0_65_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12382_ VGND VPWR VGND VPWR _07961_ _07912_ keymem.key_mem\[11\]\[24\] _07957_ _07960_
+ sky130_fd_sc_hd__a211o_2
X_24368_ VGND VPWR VPWR VGND clk _00861_ reset_n keymem.key_mem\[10\]\[105\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_69_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_129_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14121_ VPWR VGND VGND VPWR _09311_ _09399_ _09592_ _09408_ _09392_ sky130_fd_sc_hd__o22ai_2
X_23319_ VGND VPWR VGND VPWR _07199_ _03981_ _07198_ _07197_ sky130_fd_sc_hd__and3b_2
XFILLER_0_65_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24299_ VGND VPWR VPWR VGND clk _00792_ reset_n keymem.key_mem\[10\]\[36\] sky130_fd_sc_hd__dfrtp_2
X_14052_ VPWR VGND VGND VPWR _09524_ key[128] _09523_ sky130_fd_sc_hd__nand2_2
XFILLER_0_238_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13003_ VGND VPWR enc_block.round_key\[83\] _08522_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_247_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_265_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18860_ VGND VPWR VGND VPWR _04704_ _04703_ _04705_ _04077_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_101_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17811_ VGND VPWR VGND VPWR _03178_ _03792_ _03795_ _03793_ _03727_ _03803_ sky130_fd_sc_hd__a2111oi_2
X_18791_ VPWR VGND VPWR VGND _04642_ block[36] _04351_ enc_block.block_w1_reg\[4\]
+ _03954_ _04643_ sky130_fd_sc_hd__a221o_2
XFILLER_0_234_524 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_179_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17742_ VGND VPWR _00178_ _03759_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_175_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14954_ VPWR VGND VPWR VGND _10418_ enc_block.block_w0_reg\[12\] _09273_ sky130_fd_sc_hd__or2_2
XFILLER_0_27_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_136_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13905_ VPWR VGND VPWR VGND _09299_ _09317_ _09300_ _09254_ _09377_ sky130_fd_sc_hd__or4_2
XFILLER_0_175_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17673_ VGND VPWR VPWR VGND _03703_ _03711_ keymem.prev_key0_reg\[16\] _03712_ sky130_fd_sc_hd__mux2_2
X_14885_ VPWR VGND VGND VPWR _09110_ _10350_ _09097_ sky130_fd_sc_hd__nor2_2
XFILLER_0_72_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_102_1_Right_703 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_255_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19412_ VGND VPWR _05102_ _05094_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_216_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16624_ VGND VPWR VGND VPWR _02777_ _02778_ _02780_ _02776_ sky130_fd_sc_hd__nand3_2
X_13836_ VGND VPWR VGND VPWR _09308_ _09289_ _09288_ keymem.prev_key1_reg\[28\] _09003_
+ _09002_ sky130_fd_sc_hd__a32o_2
XFILLER_0_58_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19343_ VPWR VGND keymem.key_mem_we _05056_ _03560_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16555_ VPWR VGND _02714_ keymem.prev_key1_reg\[57\] keymem.prev_key1_reg\[25\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
X_13767_ VPWR VGND _09165_ _09239_ _09238_ VPWR VGND sky130_fd_sc_hd__and2_2
X_15506_ VGND VPWR VGND VPWR _10965_ _10732_ _10916_ _10963_ _10966_ sky130_fd_sc_hd__a31o_2
X_19274_ VGND VPWR _00458_ _05011_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12718_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[55\] _07651_ keymem.key_mem\[1\]\[55\]
+ _07855_ _08266_ sky130_fd_sc_hd__a22o_2
X_16486_ VGND VPWR _02647_ _09988_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13698_ VGND VPWR VGND VPWR _09170_ _09168_ _09113_ _09167_ _09067_ _09169_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_45_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_112_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_721 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_186_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18225_ VPWR VGND VPWR VGND _04133_ enc_block.round_key\[110\] _04132_ sky130_fd_sc_hd__or2_2
X_15437_ _10895_ _10898_ _10894_ _10897_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_12649_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[49\] _07744_ keymem.key_mem\[12\]\[49\]
+ _07806_ _08203_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_183_2_Right_255 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_245_1116 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_147_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_127_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18156_ _04068_ _04070_ _04065_ _04069_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_83_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_25_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15368_ VGND VPWR _10830_ keymem.prev_key1_reg\[10\] keymem.prev_key1_reg\[42\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_147_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_227_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17107_ VPWR VGND VGND VPWR _02647_ _03223_ key[68] sky130_fd_sc_hd__nor2_2
X_14319_ VPWR VGND VGND VPWR _09769_ _09779_ _09788_ _09789_ sky130_fd_sc_hd__nor3_2
XFILLER_0_83_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18087_ VPWR VGND VPWR VGND _04006_ _03992_ _04003_ enc_block.block_w0_reg\[2\] _03976_
+ _00276_ sky130_fd_sc_hd__a221o_2
X_15299_ VPWR VGND VGND VPWR _10565_ _10761_ _10480_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_307 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_1088 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17038_ VGND VPWR VGND VPWR _03161_ _03152_ key[189] _03155_ _03160_ sky130_fd_sc_hd__a211o_2
XFILLER_0_22_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1196 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18989_ VPWR VGND VGND VPWR _04778_ _04821_ _04240_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_193_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_268 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_217_1218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20951_ VGND VPWR _01224_ _05922_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_234_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_590 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_205_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23670_ keymem.prev_key0_reg\[26\] clk _00167_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_7_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20882_ VGND VPWR _01192_ _05885_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_152_1254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22621_ VGND VPWR _02036_ _06780_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_187_1306 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25340_ VGND VPWR VPWR VGND clk _01833_ reset_n keymem.key_mem\[2\]\[53\] sky130_fd_sc_hd__dfrtp_2
X_22552_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[78\] _06754_ _06753_ _04997_ _01986_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_9_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_710 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_130_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_442 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21503_ VGND VPWR _01484_ _06214_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_267_1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25271_ VGND VPWR VPWR VGND clk _01764_ reset_n keymem.key_mem\[3\]\[112\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_173_350 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_118_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22483_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[36\] _06707_ _06706_ _04927_ _01944_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_133_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_267_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24222_ VGND VPWR VPWR VGND clk _00715_ reset_n keymem.key_mem\[11\]\[87\] sky130_fd_sc_hd__dfrtp_2
X_21434_ VGND VPWR _01451_ _06178_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_71_370 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_86_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24153_ VGND VPWR VPWR VGND clk _00646_ reset_n keymem.key_mem\[11\]\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21365_ VGND VPWR _01418_ _06142_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_4_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23104_ VGND VPWR _02270_ _07029_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20316_ VGND VPWR VPWR VGND _05580_ _02998_ keymem.key_mem\[9\]\[44\] _05584_ sky130_fd_sc_hd__mux2_2
X_24084_ VGND VPWR VPWR VGND clk _00577_ reset_n keymem.key_mem\[12\]\[77\] sky130_fd_sc_hd__dfrtp_2
X_21296_ VGND VPWR _01387_ _06104_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_202_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23035_ VGND VPWR VGND VPWR _03281_ key[195] _09928_ _06987_ sky130_fd_sc_hd__a21o_2
X_20247_ VPWR VGND VGND VPWR _05548_ keymem.key_mem\[9\]\[11\] _05532_ sky130_fd_sc_hd__nand2_2
XFILLER_0_257_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20178_ VGND VPWR _00864_ _05509_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_244_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24986_ VGND VPWR VPWR VGND clk _01479_ reset_n keymem.key_mem\[5\]\[83\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_235_1318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23937_ VGND VPWR VPWR VGND clk _00430_ reset_n keymem.key_mem\[13\]\[58\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_197_910 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11951_ VGND VPWR VGND VPWR _07526_ _07554_ _07525_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_58_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14670_ VPWR VGND _09582_ _10137_ _09391_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_19_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11882_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[12\] dec_new_block\[108\]
+ _07505_ sky130_fd_sc_hd__mux2_2
X_23868_ VGND VPWR VPWR VGND clk _00361_ reset_n enc_block.block_w2_reg\[21\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_312 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13621_ VPWR VGND VPWR VGND _09092_ _09093_ _09078_ _09084_ sky130_fd_sc_hd__or3b_2
X_25607_ VGND VPWR VPWR VGND clk _02100_ reset_n keymem.key_mem\[0\]\[64\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_197_998 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_196_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22819_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[118\] _06860_ _06859_ _05071_ _02154_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_170_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23799_ VGND VPWR VPWR VGND clk _00292_ reset_n enc_block.block_w0_reg\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16340_ VPWR VGND VPWR VGND _02501_ _02502_ _02503_ _11335_ _11371_ sky130_fd_sc_hd__or4b_2
XFILLER_0_66_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13552_ VGND VPWR VGND VPWR _09024_ enc_block.block_w2_reg\[0\] enc_block.sword_ctr_reg\[1\]
+ enc_block.sword_ctr_reg\[0\] sky130_fd_sc_hd__and3b_2
XFILLER_0_251_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25538_ VGND VPWR VPWR VGND clk _02031_ reset_n keymem.key_mem\[1\]\[123\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_66_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12503_ VPWR VGND VPWR VGND keymem.key_mem\[4\]\[35\] _07734_ keymem.key_mem\[1\]\[35\]
+ _07969_ _08071_ sky130_fd_sc_hd__a22o_2
X_16271_ VPWR VGND VPWR VGND _11401_ _02434_ _11405_ _11394_ _02435_ sky130_fd_sc_hd__or4_2
X_13483_ VGND VPWR _08955_ _08954_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_246_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25469_ VGND VPWR VPWR VGND clk _01962_ reset_n keymem.key_mem\[1\]\[54\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_81_156 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18010_ VGND VPWR VGND VPWR _03736_ keymem.prev_key0_reg\[126\] _03938_ _00267_ sky130_fd_sc_hd__a21o_2
X_15222_ VGND VPWR VGND VPWR _10480_ _10602_ _10482_ _10612_ _10685_ sky130_fd_sc_hd__o22a_2
XFILLER_0_129_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12434_ VGND VPWR _08008_ _07547_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_35_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_247 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_69_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15153_ VPWR VGND VPWR VGND _10606_ _10616_ _10617_ _10589_ _10597_ sky130_fd_sc_hd__or4b_2
X_12365_ VPWR VGND VPWR VGND _07944_ keymem.key_mem\[3\]\[23\] _07619_ keymem.key_mem\[10\]\[23\]
+ _07629_ _07945_ sky130_fd_sc_hd__a221o_2
XFILLER_0_50_554 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_65_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14104_ VPWR VGND VPWR VGND _09571_ _09574_ _09572_ _09448_ _09575_ sky130_fd_sc_hd__or4_2
X_15084_ VGND VPWR VGND VPWR _10543_ _10547_ _10498_ _10536_ _10548_ sky130_fd_sc_hd__o22a_2
X_19961_ VGND VPWR _00761_ _05395_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12296_ VGND VPWR VGND VPWR _07882_ _07877_ keymem.key_mem\[10\]\[17\] _07879_ _07881_
+ sky130_fd_sc_hd__a211o_2
XPHY_EDGE_ROW_168_1_Left_435 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18912_ VPWR VGND VGND VPWR _04654_ _04752_ _04159_ sky130_fd_sc_hd__nor2_2
X_14035_ VGND VPWR VGND VPWR _09239_ keymem.round_ctr_reg\[0\] _09507_ _09506_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_129_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19892_ VGND VPWR _00730_ _05357_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_136_2_Left_607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18843_ VGND VPWR VGND VPWR _04688_ enc_block.round_key\[41\] _04149_ _04690_ sky130_fd_sc_hd__a21o_2
X_18774_ VGND VPWR _04627_ enc_block.block_w1_reg\[2\] _04626_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15986_ VPWR VGND VGND VPWR _10735_ _11161_ _11441_ _11442_ sky130_fd_sc_hd__nor3_2
XFILLER_0_234_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17725_ VPWR VGND VGND VPWR _03749_ _03750_ _03731_ sky130_fd_sc_hd__nor2_2
X_14937_ VPWR VGND VPWR VGND _10401_ enc_block.block_w0_reg\[10\] _09273_ sky130_fd_sc_hd__or2_2
XFILLER_0_76_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_76_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17656_ VGND VPWR VPWR VGND _03691_ key[139] keymem.prev_key1_reg\[11\] _03700_ sky130_fd_sc_hd__mux2_2
XFILLER_0_159_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_37_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14868_ VGND VPWR VGND VPWR _09687_ _09110_ _09146_ _09125_ _10333_ sky130_fd_sc_hd__o22a_2
XPHY_EDGE_ROW_103_1_Right_704 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_230_560 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_203_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16607_ VPWR VGND VPWR VGND _02763_ _02677_ _02754_ key[155] _02723_ _02764_ sky130_fd_sc_hd__a221o_2
X_13819_ VGND VPWR _09291_ _09290_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_230_582 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17587_ VPWR VGND VPWR VGND _03646_ _03643_ _03642_ key[252] _08929_ _03647_ sky130_fd_sc_hd__a221o_2
XFILLER_0_159_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14799_ VGND VPWR _10265_ keymem.prev_key0_reg\[38\] keymem.prev_key0_reg\[70\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_147_328 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_58_665 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19326_ VGND VPWR _00477_ _05044_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16538_ VGND VPWR VGND VPWR _11532_ _11502_ keymem.rcon_logic.tmp_rcon\[2\] _02697_
+ sky130_fd_sc_hd__a21o_2
XFILLER_0_45_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_57_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_162_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19257_ VPWR VGND keymem.key_mem\[13\]\[80\] _05001_ _04979_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16469_ VGND VPWR VGND VPWR _02629_ _02628_ _02630_ _02627_ _02626_ sky130_fd_sc_hd__nand4_2
X_18208_ VPWR VGND VPWR VGND _04117_ _04040_ _04115_ enc_block.block_w0_reg\[12\]
+ _04097_ _00286_ sky130_fd_sc_hd__a221o_2
XFILLER_0_115_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_434 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_562 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_147_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19188_ VGND VPWR _00424_ _04959_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_184_2_Right_256 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_83_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18139_ VGND VPWR _04054_ enc_block.block_w2_reg\[15\] enc_block.block_w1_reg\[23\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1391 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_48_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21150_ VGND VPWR VPWR VGND _06018_ _03056_ keymem.key_mem\[6\]\[50\] _06028_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_68_2_Left_539 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_651 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20101_ VGND VPWR _05469_ _05387_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21081_ VGND VPWR VPWR VGND _05983_ _11546_ keymem.key_mem\[6\]\[17\] _05992_ sky130_fd_sc_hd__mux2_2
X_20032_ VGND VPWR VPWR VGND _05424_ _02945_ keymem.key_mem\[10\]\[39\] _05433_ sky130_fd_sc_hd__mux2_2
XFILLER_0_119_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24840_ VGND VPWR VPWR VGND clk _01333_ reset_n keymem.key_mem\[6\]\[65\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21983_ VGND VPWR _01707_ _06471_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24771_ VGND VPWR VPWR VGND clk _01264_ reset_n keymem.key_mem\[7\]\[124\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_55_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23722_ keymem.prev_key0_reg\[78\] clk _00219_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20934_ VGND VPWR _01216_ _05913_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_55_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_182_2_Left_653 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_234_1373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20865_ VGND VPWR _01184_ _05876_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23653_ keymem.prev_key0_reg\[9\] clk _00150_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_138_339 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22604_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[114\] _06777_ _06776_ _05062_ _02022_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_37_827 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_64_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23584_ VGND VPWR VPWR VGND clk _00085_ reset_n keymem.key_mem\[14\]\[73\] sky130_fd_sc_hd__dfrtp_2
X_20796_ VGND VPWR VGND VPWR _05839_ keymem.key_mem_we _10977_ _05838_ _01152_ sky130_fd_sc_hd__a31o_2
XFILLER_0_48_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22535_ VGND VPWR _01975_ _06755_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25323_ VGND VPWR VPWR VGND clk _01816_ reset_n keymem.key_mem\[2\]\[36\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_64_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_10_1029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_819 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_221_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_228_1122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_49_1228 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_267_1182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25254_ VGND VPWR VPWR VGND clk _01747_ reset_n keymem.key_mem\[3\]\[95\] sky130_fd_sc_hd__dfrtp_2
X_22466_ VGND VPWR _01934_ _06727_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_63_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_66_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21417_ VGND VPWR _01443_ _06169_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24205_ VGND VPWR VPWR VGND clk _00698_ reset_n keymem.key_mem\[11\]\[70\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_543 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25185_ VGND VPWR VPWR VGND clk _01678_ reset_n keymem.key_mem\[3\]\[26\] sky130_fd_sc_hd__dfrtp_2
X_22397_ VGND VPWR VPWR VGND _06680_ _03640_ keymem.key_mem\[2\]\[123\] _06690_ sky130_fd_sc_hd__mux2_2
XFILLER_0_161_386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_874 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_716 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_280 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12150_ VGND VPWR _07746_ _07571_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24136_ VGND VPWR VPWR VGND clk _00629_ reset_n keymem.key_mem\[11\]\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_206_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21348_ VGND VPWR _01410_ _06133_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_202_1317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24067_ VGND VPWR VPWR VGND clk _00560_ reset_n keymem.key_mem\[12\]\[60\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_206_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12081_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[4\] _07585_ keymem.key_mem\[7\]\[4\]
+ _07566_ _07680_ sky130_fd_sc_hd__a22o_2
X_21279_ VGND VPWR _01379_ _06095_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23018_ VGND VPWR VGND VPWR _03133_ _06928_ _03138_ _06978_ sky130_fd_sc_hd__a21o_2
XFILLER_0_200_1030 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_263_438 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_102_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1196 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_228_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15840_ VGND VPWR _11296_ _11295_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_137_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_825 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_176_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15771_ VGND VPWR _11227_ _11192_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24969_ VGND VPWR VPWR VGND clk _01462_ reset_n keymem.key_mem\[5\]\[66\] sky130_fd_sc_hd__dfrtp_2
X_12983_ VGND VPWR enc_block.round_key\[81\] _08504_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_137_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1070 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17510_ VPWR VGND VPWR VGND _03579_ _03494_ _03575_ key[242] _03527_ _03580_ sky130_fd_sc_hd__a221o_2
XFILLER_0_73_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14722_ VGND VPWR _10189_ _09987_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18490_ VGND VPWR _04372_ enc_block.block_w3_reg\[14\] enc_block.block_w2_reg\[22\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_11934_ VGND VPWR VGND VPWR _07529_ _07537_ _07528_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_891 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_212_582 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17441_ VPWR VGND VGND VPWR _03520_ _03240_ _02957_ sky130_fd_sc_hd__nand2_2
X_14653_ VPWR VGND VPWR VGND _10112_ _10119_ _10117_ _10110_ _10120_ sky130_fd_sc_hd__or4_2
XFILLER_0_196_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_213_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11865_ VGND VPWR result[99] _07496_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_39_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13604_ VPWR VGND VPWR VGND _09013_ _08997_ _09034_ _09001_ _09076_ sky130_fd_sc_hd__or4_2
XFILLER_0_131_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17372_ VGND VPWR VPWR VGND _03384_ keymem.key_mem\[14\]\[95\] _03460_ _03461_ sky130_fd_sc_hd__mux2_2
X_14584_ VPWR VGND VGND VPWR _09408_ _10052_ _09294_ sky130_fd_sc_hd__nor2_2
XFILLER_0_28_838 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11796_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[1\] dec_new_block\[65\]
+ _07462_ sky130_fd_sc_hd__mux2_2
XFILLER_0_248_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_158 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19111_ VPWR VGND keymem.key_mem\[13\]\[24\] _04911_ _04903_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16323_ VGND VPWR _02485_ _10993_ _02486_ _11018_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_13535_ VGND VPWR _09007_ _09006_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_55_657 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_55_679 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_137_383 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19042_ VPWR VGND VPWR VGND _04867_ _04788_ _04866_ enc_block.block_w2_reg\[30\]
+ _04613_ _00370_ sky130_fd_sc_hd__a221o_2
XFILLER_0_10_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16254_ VGND VPWR _11338_ _11211_ _02418_ _11280_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_42_329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13466_ VGND VPWR VGND VPWR aes_core_ctrl_reg\[0\] init aes_core_ctrl_reg\[2\] _08938_
+ sky130_fd_sc_hd__a21o_2
XFILLER_0_35_370 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15205_ VGND VPWR _10668_ _10496_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_51_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12417_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[27\] _07644_ _07992_ _07988_ _07993_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_3_949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16185_ VGND VPWR VGND VPWR _02350_ _02345_ _11338_ _02347_ _02349_ sky130_fd_sc_hd__a211o_2
X_13397_ VGND VPWR VGND VPWR _08877_ _07579_ keymem.key_mem\[12\]\[123\] _08876_ _07616_
+ sky130_fd_sc_hd__a211o_2
X_15136_ VPWR VGND VGND VPWR _10583_ _10600_ _10496_ sky130_fd_sc_hd__nor2_2
XFILLER_0_267_722 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_236_Right_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_224_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12348_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[21\] _07683_ keymem.key_mem\[8\]\[21\]
+ _07929_ _07930_ sky130_fd_sc_hd__a22o_2
XFILLER_0_11_749 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15067_ VGND VPWR VGND VPWR _10459_ _10527_ _10528_ _10530_ _10531_ sky130_fd_sc_hd__a31o_2
X_12279_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[16\] _07865_ keymem.key_mem\[12\]\[16\]
+ _07621_ _07866_ sky130_fd_sc_hd__a22o_2
X_19944_ VGND VPWR _00755_ _05384_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_267_788 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_142_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14018_ VGND VPWR VPWR VGND _09489_ _09431_ _09426_ _09490_ sky130_fd_sc_hd__or3_2
X_19875_ VGND VPWR _00722_ _05348_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18826_ VPWR VGND VPWR VGND _04674_ _04664_ _04673_ enc_block.block_w2_reg\[7\] _04602_
+ _00347_ sky130_fd_sc_hd__a221o_2
XFILLER_0_250_600 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_223_836 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18757_ VPWR VGND _04612_ _04611_ enc_block.round_key\[33\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15969_ VPWR VGND VGND VPWR _11245_ _11326_ _11425_ _11385_ _11370_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_218_1368 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17708_ VGND VPWR _03738_ _03281_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_218_1379 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18688_ VGND VPWR _04550_ _03949_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_231_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17639_ VGND VPWR _00146_ _03688_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_104_1_Right_705 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20650_ VGND VPWR VGND VPWR _05676_ _03279_ _01086_ _05759_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_110_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_85_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19309_ VPWR VGND keymem.key_mem_we _05033_ _03492_ VPWR VGND sky130_fd_sc_hd__and2_2
X_20581_ VGND VPWR _01053_ _05723_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_2_1141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_721 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22320_ VGND VPWR VPWR VGND _06647_ _03383_ keymem.key_mem\[2\]\[86\] _06650_ sky130_fd_sc_hd__mux2_2
XFILLER_0_2_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_143_364 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22251_ VGND VPWR VPWR VGND _06611_ _03082_ keymem.key_mem\[2\]\[53\] _06614_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_185_2_Right_257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_170_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21202_ VGND VPWR _06055_ _03279_ _01342_ _05985_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_223_1030 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22182_ VGND VPWR _01800_ _06577_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_160_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21133_ VGND VPWR _01309_ _06019_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_2_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_121_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21064_ VGND VPWR _01277_ _05982_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_226_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20015_ VGND VPWR _05424_ _05388_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_119_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24823_ VGND VPWR VPWR VGND clk _01316_ reset_n keymem.key_mem\[6\]\[48\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24754_ VGND VPWR VPWR VGND clk _01247_ reset_n keymem.key_mem\[7\]\[107\] sky130_fd_sc_hd__dfrtp_2
X_21966_ VGND VPWR _06462_ _06402_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_16_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23705_ keymem.prev_key0_reg\[61\] clk _00202_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20917_ VGND VPWR VPWR VGND _01208_ _05824_ _03226_ _08922_ _05904_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_171_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24685_ VGND VPWR VPWR VGND clk _01178_ reset_n keymem.key_mem\[7\]\[38\] sky130_fd_sc_hd__dfrtp_2
X_21897_ VPWR VGND keymem.key_mem\[3\]\[16\] _06425_ _06413_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_51_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11650_ VGND VPWR _07387_ _07386_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20848_ VGND VPWR VPWR VGND _05867_ _04927_ keymem.key_mem\[7\]\[36\] _05868_ sky130_fd_sc_hd__mux2_2
X_23636_ VGND VPWR VPWR VGND clk _00137_ reset_n keymem.key_mem\[14\]\[125\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_484 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_36_112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23567_ VGND VPWR VPWR VGND clk _00068_ reset_n keymem.key_mem\[14\]\[56\] sky130_fd_sc_hd__dfrtp_2
X_20779_ VGND VPWR _05830_ _05823_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25306_ VGND VPWR VPWR VGND clk _01799_ reset_n keymem.key_mem\[2\]\[19\] sky130_fd_sc_hd__dfrtp_2
X_13320_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[115\] _07748_ keymem.key_mem\[12\]\[115\]
+ _07722_ _08808_ sky130_fd_sc_hd__a22o_2
X_22518_ VGND VPWR _01967_ _06746_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23498_ VPWR VGND VGND VPWR _07358_ _07167_ _07357_ sky130_fd_sc_hd__nand2_2
XFILLER_0_165_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25237_ VGND VPWR VPWR VGND clk _01730_ reset_n keymem.key_mem\[3\]\[78\] sky130_fd_sc_hd__dfrtp_2
X_22449_ VGND VPWR _01926_ _06718_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13251_ VGND VPWR VGND VPWR _07542_ keymem.key_mem\[8\]\[108\] _08743_ _08745_ _08746_
+ _08736_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_27_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12202_ VGND VPWR enc_block.round_key\[10\] _07794_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13182_ VPWR VGND VPWR VGND _08683_ keymem.key_mem\[13\]\[101\] _08125_ keymem.key_mem\[9\]\[101\]
+ _07919_ _08684_ sky130_fd_sc_hd__a221o_2
XFILLER_0_27_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_682 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25168_ VGND VPWR VPWR VGND clk _01661_ reset_n keymem.key_mem\[3\]\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_206_1261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12133_ VGND VPWR enc_block.round_key\[6\] _07729_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24119_ VGND VPWR VPWR VGND clk _00612_ reset_n keymem.key_mem\[12\]\[112\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_102_272 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25099_ VGND VPWR VPWR VGND clk _01592_ reset_n keymem.key_mem\[4\]\[68\] sky130_fd_sc_hd__dfrtp_2
X_17990_ VGND VPWR VGND VPWR _02647_ keymem.prev_key1_reg\[120\] _03679_ _03925_ sky130_fd_sc_hd__a21o_2
XFILLER_0_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16941_ VPWR VGND VPWR VGND keymem.prev_key1_reg\[52\] _03073_ _02473_ _02474_ sky130_fd_sc_hd__or3b_2
X_12064_ VGND VPWR VGND VPWR _07648_ keymem.key_mem\[2\]\[3\] _07653_ _07661_ _07664_
+ _07663_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_236_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_198_1062 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19660_ VGND VPWR VPWR VGND _05227_ _05079_ keymem.key_mem\[12\]\[122\] _05234_ sky130_fd_sc_hd__mux2_2
XFILLER_0_99_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16872_ VGND VPWR VGND VPWR _03009_ _09796_ _11055_ _11092_ _03010_ sky130_fd_sc_hd__a31o_2
X_18611_ VGND VPWR _04481_ enc_block.block_w3_reg\[9\] enc_block.block_w3_reg\[10\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15823_ VGND VPWR VPWR VGND _11265_ _11247_ _11233_ _11279_ sky130_fd_sc_hd__or3_2
XFILLER_0_137_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19591_ VGND VPWR VPWR VGND _05183_ _05015_ keymem.key_mem\[12\]\[89\] _05198_ sky130_fd_sc_hd__mux2_2
X_18542_ VPWR VGND VGND VPWR _04419_ _04343_ _04417_ sky130_fd_sc_hd__nand2_2
XFILLER_0_99_362 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_666 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15754_ VGND VPWR _11210_ _11209_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12966_ VPWR VGND VPWR VGND _08488_ keymem.key_mem\[13\]\[80\] _07694_ keymem.key_mem\[2\]\[80\]
+ _07646_ _08489_ sky130_fd_sc_hd__a221o_2
XFILLER_0_176_209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14705_ VPWR VGND VPWR VGND _10170_ _10171_ _10172_ _10169_ _09998_ sky130_fd_sc_hd__or4b_2
X_11917_ VGND VPWR result[125] _07522_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18473_ VPWR VGND VPWR VGND _04357_ _04353_ _04356_ sky130_fd_sc_hd__or2_2
X_15685_ VPWR VGND VGND VPWR _11142_ _11113_ _11141_ sky130_fd_sc_hd__nand2_2
X_12897_ VGND VPWR VGND VPWR _08427_ _07902_ keymem.key_mem\[11\]\[73\] _08426_ _07572_
+ sky130_fd_sc_hd__a211o_2
X_17424_ VPWR VGND VPWR VGND _03505_ _03494_ _03502_ key[230] _03366_ _03506_ sky130_fd_sc_hd__a221o_2
XFILLER_0_150_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14636_ VGND VPWR VPWR VGND _09730_ _10101_ key[133] _10103_ sky130_fd_sc_hd__mux2_2
X_11848_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[27\] dec_new_block\[91\]
+ _07488_ sky130_fd_sc_hd__mux2_2
XFILLER_0_67_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17355_ VGND VPWR _00105_ _03445_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14567_ VGND VPWR VGND VPWR _09358_ _09381_ _09355_ _09419_ _10035_ sky130_fd_sc_hd__o22a_2
X_11779_ VGND VPWR result[56] _07453_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_184_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16306_ VGND VPWR VGND VPWR _10960_ keymem.prev_key1_reg\[116\] _02470_ _10948_ sky130_fd_sc_hd__nand3_2
XFILLER_0_27_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13518_ VGND VPWR VGND VPWR _08990_ _08988_ _08987_ keymem.prev_key1_reg\[5\] _08989_
+ _08983_ sky130_fd_sc_hd__a32o_2
X_17286_ VGND VPWR _03384_ _09540_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14498_ VGND VPWR _09106_ _09219_ _09967_ _09012_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_148_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19025_ VPWR VGND VGND VPWR _04778_ _04853_ _04274_ sky130_fd_sc_hd__nor2_2
X_16237_ VGND VPWR _02402_ keymem.prev_key1_reg\[115\] _02344_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_13449_ VPWR VGND VPWR VGND _08923_ enc_block.sword_ctr_inc sky130_fd_sc_hd__inv_2
XFILLER_0_45_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_885 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_23_362 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16168_ VGND VPWR _11622_ keymem.prev_key0_reg\[114\] _11621_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_140_356 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_109_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15119_ VGND VPWR _10583_ _10502_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_107_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16099_ VGND VPWR VGND VPWR _10814_ _10775_ keymem.prev_key1_reg\[114\] _11553_ sky130_fd_sc_hd__a21o_2
XFILLER_0_259_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_220_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19927_ VGND VPWR VPWR VGND _05372_ keymem.key_mem\[11\]\[119\] _03613_ _05376_ sky130_fd_sc_hd__mux2_2
XFILLER_0_259_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19858_ VGND VPWR VPWR VGND _05339_ keymem.key_mem\[11\]\[86\] _03383_ _05340_ sky130_fd_sc_hd__mux2_2
XFILLER_0_177_1157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18809_ VPWR VGND VPWR VGND _04659_ _04656_ _04658_ sky130_fd_sc_hd__or2_2
X_19789_ VGND VPWR VPWR VGND _05303_ keymem.key_mem\[11\]\[53\] _03083_ _05304_ sky130_fd_sc_hd__mux2_2
X_21820_ VGND VPWR VPWR VGND _06377_ _03555_ keymem.key_mem\[4\]\[110\] _06382_ sky130_fd_sc_hd__mux2_2
XFILLER_0_56_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21751_ VGND VPWR VPWR VGND _06344_ _03306_ keymem.key_mem\[4\]\[77\] _06346_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20702_ VGND VPWR VPWR VGND _05783_ _03485_ keymem.key_mem\[8\]\[99\] _05787_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_105_1_Right_706 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21682_ VGND VPWR VPWR VGND _06308_ _02998_ keymem.key_mem\[4\]\[44\] _06310_ sky130_fd_sc_hd__mux2_2
X_24470_ VGND VPWR VPWR VGND clk _00963_ reset_n keymem.key_mem\[9\]\[79\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_108_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23421_ VGND VPWR _07290_ _04211_ _02326_ _07096_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_20633_ VGND VPWR VPWR VGND _05747_ _03209_ keymem.key_mem\[8\]\[66\] _05751_ sky130_fd_sc_hd__mux2_2
XFILLER_0_11_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23352_ VPWR VGND VPWR VGND _07229_ enc_block.round_key\[14\] _07227_ sky130_fd_sc_hd__or2_2
XFILLER_0_11_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20564_ VGND VPWR VPWR VGND _05714_ _02883_ keymem.key_mem\[8\]\[33\] _05715_ sky130_fd_sc_hd__mux2_2
XFILLER_0_6_562 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22303_ VGND VPWR VPWR VGND _06634_ _03314_ keymem.key_mem\[2\]\[78\] _06641_ sky130_fd_sc_hd__mux2_2
XFILLER_0_150_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23283_ VPWR VGND _07166_ enc_block.block_w2_reg\[0\] enc_block.block_w3_reg\[24\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_225_1114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_131_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20495_ VGND VPWR VPWR VGND _05676_ _09724_ keymem.key_mem\[8\]\[1\] _05678_ sky130_fd_sc_hd__mux2_2
XFILLER_0_127_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22234_ VGND VPWR VPWR VGND _06600_ _03006_ keymem.key_mem\[2\]\[45\] _06605_ sky130_fd_sc_hd__mux2_2
X_25022_ VGND VPWR VPWR VGND clk _01515_ reset_n keymem.key_mem\[5\]\[119\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_186_2_Right_258 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_258_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22165_ VGND VPWR VPWR VGND _06565_ _10976_ keymem.key_mem\[2\]\[12\] _06569_ sky130_fd_sc_hd__mux2_2
XFILLER_0_203_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21116_ VGND VPWR _01301_ _06010_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_160_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22096_ VGND VPWR VPWR VGND _06527_ _05052_ keymem.key_mem\[3\]\[109\] _06531_ sky130_fd_sc_hd__mux2_2
XFILLER_0_246_769 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_22_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_227_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21047_ VGND VPWR VPWR VGND _05972_ _09724_ keymem.key_mem\[6\]\[1\] _05974_ sky130_fd_sc_hd__mux2_2
XFILLER_0_226_460 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_156_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_835 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_260_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_96_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_242_975 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_241_Left_508 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12820_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[65\] _08259_ _08357_ _08353_ _08358_
+ sky130_fd_sc_hd__o22a_2
X_24806_ VGND VPWR VPWR VGND clk _01299_ reset_n keymem.key_mem\[6\]\[31\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_198_345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25786_ keymem.prev_key1_reg\[102\] clk _02279_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22998_ VPWR VGND VPWR VGND _06966_ _03066_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_485 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12751_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[58\] _07793_ _08295_ _08291_ _08296_
+ sky130_fd_sc_hd__o22a_2
X_24737_ VGND VPWR VPWR VGND clk _01230_ reset_n keymem.key_mem\[7\]\[90\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_214_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21949_ VGND VPWR _01691_ _06453_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_96_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11702_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[18\] dec_new_block\[18\]
+ _07415_ sky130_fd_sc_hd__mux2_2
X_15470_ VPWR VGND VPWR VGND _10925_ _10929_ _10926_ _10438_ _10930_ sky130_fd_sc_hd__or4_2
XFILLER_0_132_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12682_ VPWR VGND VPWR VGND _08232_ keymem.key_mem\[14\]\[52\] _08003_ keymem.key_mem\[12\]\[52\]
+ _07807_ _08233_ sky130_fd_sc_hd__a221o_2
X_24668_ VGND VPWR VPWR VGND clk _01161_ reset_n keymem.key_mem\[7\]\[21\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_177_1_Left_444 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_166_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14421_ VGND VPWR VGND VPWR _09466_ _09355_ _09476_ _09890_ sky130_fd_sc_hd__a21o_2
X_11633_ VPWR VGND VPWR VGND _07373_ enc_block.enc_ctrl_reg\[3\] enc_block.enc_ctrl_reg\[2\]
+ sky130_fd_sc_hd__or2_2
X_23619_ VGND VPWR VPWR VGND clk _00120_ reset_n keymem.key_mem\[14\]\[108\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_145_2_Left_616 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_112_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24599_ VGND VPWR VPWR VGND clk _01092_ reset_n keymem.key_mem\[8\]\[80\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17140_ VGND VPWR VPWR VGND _03185_ keymem.key_mem\[14\]\[71\] _03252_ _03253_ sky130_fd_sc_hd__mux2_2
X_14352_ VGND VPWR _09821_ _09106_ _09822_ _09818_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_52_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_167_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_958 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_247_1361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_250_Left_517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13303_ VGND VPWR VGND VPWR _08793_ _07968_ keymem.key_mem\[9\]\[113\] _08790_ _08792_
+ sky130_fd_sc_hd__a211o_2
X_17071_ VPWR VGND VPWR VGND _03191_ keymem.prev_key0_reg\[64\] _09717_ _09508_ _09721_
+ _03190_ sky130_fd_sc_hd__o311a_2
X_14283_ VGND VPWR VGND VPWR _09399_ _09456_ _09330_ _09441_ _09753_ sky130_fd_sc_hd__o22a_2
XFILLER_0_40_608 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_243_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16022_ VGND VPWR _11477_ _11247_ _11221_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_13234_ VGND VPWR VGND VPWR _08731_ _07721_ keymem.key_mem\[14\]\[106\] _08728_ _08730_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_27_1142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_855 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13165_ VGND VPWR enc_block.round_key\[99\] _08668_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_236_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12116_ VPWR VGND VPWR VGND keymem.key_mem\[4\]\[6\] _07693_ keymem.key_mem\[2\]\[6\]
+ _07647_ _07713_ sky130_fd_sc_hd__a22o_2
X_17973_ VGND VPWR VPWR VGND _03896_ _03913_ keymem.prev_key0_reg\[114\] _03914_ sky130_fd_sc_hd__mux2_2
XFILLER_0_264_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13096_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[93\] _07779_ keymem.key_mem\[10\]\[93\]
+ _07785_ _08606_ sky130_fd_sc_hd__a22o_2
XFILLER_0_209_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_100_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_137_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16924_ VGND VPWR _00062_ _03057_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19712_ VGND VPWR _00644_ _05263_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12047_ VGND VPWR _07647_ _07646_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_137_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_40_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16855_ VPWR VGND VGND VPWR _02995_ _09732_ _10968_ sky130_fd_sc_hd__nand2_2
XFILLER_0_205_633 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19643_ VGND VPWR VPWR VGND _05216_ _05062_ keymem.key_mem\[12\]\[114\] _05225_ sky130_fd_sc_hd__mux2_2
XFILLER_0_178_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_148_2_Right_220 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15806_ VGND VPWR _11262_ _11261_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19574_ VGND VPWR VGND VPWR _05189_ keymem.key_mem_we _03330_ _05187_ _00580_ sky130_fd_sc_hd__a31o_2
XFILLER_0_254_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_217_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16786_ VGND VPWR VGND VPWR _10276_ _10275_ _02931_ _02932_ sky130_fd_sc_hd__a21o_2
XFILLER_0_254_1376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13998_ VPWR VGND VPWR VGND _09469_ _09470_ _09465_ _09467_ sky130_fd_sc_hd__or3b_2
X_18525_ VPWR VGND VGND VPWR _04403_ _04404_ _04077_ sky130_fd_sc_hd__nor2_2
X_15737_ enc_block.sword_ctr_reg\[1\] _11193_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[20\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_12949_ VGND VPWR VGND VPWR _08474_ _07593_ keymem.key_mem\[9\]\[78\] _08473_ _07616_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_141_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18456_ VGND VPWR _04341_ enc_block.block_w3_reg\[11\] _04340_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_239_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15668_ VGND VPWR VGND VPWR _11125_ _11124_ _11123_ _11122_ _11121_ sky130_fd_sc_hd__and4_2
XFILLER_0_29_933 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_77_2_Left_548 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_111_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_150_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17407_ VPWR VGND VGND VPWR _03491_ key[228] _10838_ sky130_fd_sc_hd__nand2_2
X_14619_ VPWR VGND _10056_ _10087_ _10075_ VPWR VGND sky130_fd_sc_hd__and2_2
X_18387_ _04278_ _04280_ _04008_ _04279_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_111_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_240 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15599_ VPWR VGND VGND VPWR _11057_ _10215_ _10229_ sky130_fd_sc_hd__nand2_2
XFILLER_0_28_465 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_51_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17338_ VGND VPWR _09988_ keymem.prev_key0_reg\[92\] _03430_ _02771_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_12_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_185_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_261_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17269_ VGND VPWR keymem.prev_key0_reg\[85\] _02539_ _03368_ _02540_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_24_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19008_ VGND VPWR _04837_ _03957_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_70_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_259_327 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_178_11 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_11_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20280_ VGND VPWR VPWR VGND _05558_ _02765_ keymem.key_mem\[9\]\[27\] _05565_ sky130_fd_sc_hd__mux2_2
XFILLER_0_144_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_844 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_261_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_191_2_Left_662 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_140_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_122_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_46_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23970_ VGND VPWR VPWR VGND clk _00463_ reset_n keymem.key_mem\[13\]\[91\] sky130_fd_sc_hd__dfrtp_2
X_22921_ VGND VPWR VGND VPWR _02198_ _06918_ _06916_ keymem.prev_key1_reg\[21\] sky130_fd_sc_hd__o21a_2
XFILLER_0_93_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25640_ VGND VPWR VPWR VGND clk _02133_ reset_n keymem.key_mem\[0\]\[97\] sky130_fd_sc_hd__dfrtp_2
X_22852_ VPWR VGND VPWR VGND _06874_ keymem.round_ctr_reg\[2\] _05241_ sky130_fd_sc_hd__or2_2
XFILLER_0_233_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21803_ VGND VPWR VPWR VGND _06366_ _03506_ keymem.key_mem\[4\]\[102\] _06373_ sky130_fd_sc_hd__mux2_2
XFILLER_0_190_1165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25571_ VGND VPWR VPWR VGND clk _02064_ reset_n keymem.key_mem\[0\]\[28\] sky130_fd_sc_hd__dfrtp_2
X_22783_ VGND VPWR _02126_ _06852_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24522_ VGND VPWR VPWR VGND clk _01015_ reset_n keymem.key_mem\[8\]\[3\] sky130_fd_sc_hd__dfrtp_2
X_21734_ VGND VPWR VPWR VGND _06330_ _03234_ keymem.key_mem\[4\]\[69\] _06337_ sky130_fd_sc_hd__mux2_2
XFILLER_0_133_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_106_1_Right_707 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24453_ VGND VPWR VPWR VGND clk _00946_ reset_n keymem.key_mem\[9\]\[62\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_110_2_Right_182 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21665_ VGND VPWR VPWR VGND _06297_ _02913_ keymem.key_mem\[4\]\[36\] _06301_ sky130_fd_sc_hd__mux2_2
XFILLER_0_30_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23404_ VGND VPWR _07275_ enc_block.block_w3_reg\[28\] _07274_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20616_ VGND VPWR VPWR VGND _05736_ _03129_ keymem.key_mem\[8\]\[58\] _05742_ sky130_fd_sc_hd__mux2_2
XFILLER_0_30_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_35_947 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24384_ VGND VPWR VPWR VGND clk _00877_ reset_n keymem.key_mem\[10\]\[121\] sky130_fd_sc_hd__dfrtp_2
X_21596_ VGND VPWR VPWR VGND _06263_ _09991_ keymem.key_mem\[4\]\[3\] _06265_ sky130_fd_sc_hd__mux2_2
XFILLER_0_61_243 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23335_ VPWR VGND VGND VPWR _07213_ enc_block.block_w2_reg\[4\] enc_block.block_w2_reg\[5\]
+ sky130_fd_sc_hd__nand2_2
X_20547_ VGND VPWR VPWR VGND _05703_ _02720_ keymem.key_mem\[8\]\[25\] _05706_ sky130_fd_sc_hd__mux2_2
XFILLER_0_43_980 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23266_ VPWR VGND VPWR VGND _07151_ _07148_ _07150_ sky130_fd_sc_hd__or2_2
X_20478_ VGND VPWR _01005_ _05668_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25005_ VGND VPWR VPWR VGND clk _01498_ reset_n keymem.key_mem\[5\]\[102\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_187_2_Right_259 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22217_ VGND VPWR VPWR VGND _06589_ _02923_ keymem.key_mem\[2\]\[37\] _06596_ sky130_fd_sc_hd__mux2_2
X_23197_ VGND VPWR _07088_ _07085_ _07087_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_22148_ VGND VPWR _01784_ _06559_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_140_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14970_ VPWR VGND VPWR VGND _10434_ enc_block.block_w0_reg\[15\] _08995_ sky130_fd_sc_hd__or2_2
X_22079_ VGND VPWR VPWR VGND _06516_ _05035_ keymem.key_mem\[3\]\[101\] _06522_ sky130_fd_sc_hd__mux2_2
XFILLER_0_22_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_514 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13921_ VGND VPWR VGND VPWR _09392_ _09386_ _09388_ _09389_ _09393_ sky130_fd_sc_hd__a31o_2
XFILLER_0_233_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_226_290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_251_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16640_ VGND VPWR _02795_ keymem.prev_key0_reg\[29\] _02794_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_13852_ VGND VPWR VGND VPWR _09320_ _09318_ _09324_ _09323_ sky130_fd_sc_hd__a21oi_2
X_25838_ VGND VPWR VPWR VGND clk _02331_ reset_n enc_block.block_w3_reg\[26\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_96_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_304 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12803_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[64\] _07908_ keymem.key_mem\[10\]\[64\]
+ _07786_ _08342_ sky130_fd_sc_hd__a22o_2
XFILLER_0_251_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16571_ VGND VPWR _02729_ keymem.prev_key0_reg\[58\] keymem.prev_key0_reg\[90\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
X_13783_ VGND VPWR _09255_ _08941_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25769_ keymem.prev_key1_reg\[85\] clk _02262_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_57_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18310_ VGND VPWR VGND VPWR _02536_ _11301_ _04073_ _04211_ sky130_fd_sc_hd__a21o_2
X_15522_ VPWR VGND VGND VPWR _10981_ _10514_ _10500_ sky130_fd_sc_hd__nand2_2
X_19290_ VGND VPWR VGND VPWR _05020_ keymem.key_mem_we _03444_ _04999_ _00465_ sky130_fd_sc_hd__a31o_2
X_12734_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[57\] _07809_ keymem.key_mem\[12\]\[57\]
+ _07807_ _08280_ sky130_fd_sc_hd__a22o_2
XFILLER_0_32_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18241_ VGND VPWR VGND VPWR _07374_ _07381_ _04148_ _03952_ sky130_fd_sc_hd__a21oi_2
X_15453_ VPWR VGND VGND VPWR _10914_ keymem.key_mem\[14\]\[11\] _09541_ sky130_fd_sc_hd__nand2_2
X_12665_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[50\] _07565_ keymem.key_mem\[1\]\[50\]
+ _07855_ _08218_ sky130_fd_sc_hd__a22o_2
XFILLER_0_37_251 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14404_ VGND VPWR VGND VPWR _09873_ _09353_ _09463_ _09331_ sky130_fd_sc_hd__o21a_2
X_18172_ VPWR VGND VGND VPWR _04085_ _10677_ _10728_ sky130_fd_sc_hd__nand2_2
X_15384_ VGND VPWR VGND VPWR _10628_ _10569_ _10477_ _10508_ _10845_ sky130_fd_sc_hd__o22a_2
XFILLER_0_203_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12596_ VGND VPWR enc_block.round_key\[43\] _08155_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_167_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17123_ VPWR VGND VPWR VGND _03237_ keymem.prev_key0_reg\[70\] sky130_fd_sc_hd__inv_2
XFILLER_0_0_1453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14335_ VGND VPWR VGND VPWR _09805_ _09051_ _09804_ _09803_ sky130_fd_sc_hd__o21a_2
XFILLER_0_13_608 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_68_1264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_194 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17054_ VPWR VGND _03175_ _02848_ _02847_ VPWR VGND sky130_fd_sc_hd__xor2_2
X_14266_ VPWR VGND VGND VPWR _09327_ _09350_ _09736_ _09564_ _09355_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_64_1139 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_180_1334 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_122_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1186 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16005_ VGND VPWR _11460_ _11459_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13217_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[105\] _07834_ keymem.key_mem\[8\]\[105\]
+ _08211_ _08715_ sky130_fd_sc_hd__a22o_2
X_14197_ VPWR VGND VGND VPWR _09665_ _09057_ _09174_ _09090_ _09668_ _09667_ sky130_fd_sc_hd__o221a_2
XFILLER_0_0_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13148_ VPWR VGND VPWR VGND _08652_ keymem.key_mem\[5\]\[98\] _07811_ keymem.key_mem\[10\]\[98\]
+ _07865_ _08653_ sky130_fd_sc_hd__a221o_2
XFILLER_0_249_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17956_ VGND VPWR VPWR VGND _03876_ key[237] keymem.prev_key1_reg\[109\] _03902_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_104_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13079_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[91\] _07668_ keymem.key_mem\[6\]\[91\]
+ _07818_ _08591_ sky130_fd_sc_hd__a22o_2
XFILLER_0_189_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16907_ VPWR VGND VGND VPWR _03042_ _03040_ _03041_ sky130_fd_sc_hd__nand2_2
X_17887_ VGND VPWR VPWR VGND _03812_ key[215] keymem.prev_key1_reg\[87\] _03855_ sky130_fd_sc_hd__mux2_2
XFILLER_0_178_1296 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_139_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_75_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19626_ VGND VPWR _05216_ _05091_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_79_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16838_ VPWR VGND _09730_ _02979_ _02978_ VPWR VGND sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_149_2_Right_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_215_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_164_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_580 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_156_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_75_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16769_ VPWR VGND VPWR VGND _02916_ _02915_ sky130_fd_sc_hd__inv_2
X_19557_ VPWR VGND keymem.key_mem\[12\]\[73\] _05180_ _05173_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_250_1037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_87_140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_250_1059 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18508_ VPWR VGND VGND VPWR _04388_ _04389_ enc_block.round_key\[71\] sky130_fd_sc_hd__nor2_2
XFILLER_0_75_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19488_ VGND VPWR _00540_ _05143_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_75_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18439_ VPWR VGND VPWR VGND _04325_ block[65] _04213_ enc_block.block_w0_reg\[1\]
+ _04276_ _04326_ sky130_fd_sc_hd__a221o_2
XFILLER_0_75_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_189_1370 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_12_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21450_ VGND VPWR VPWR VGND _06184_ _03183_ keymem.key_mem\[5\]\[63\] _06187_ sky130_fd_sc_hd__mux2_2
XFILLER_0_43_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_111_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20401_ VGND VPWR _00968_ _05628_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_160_215 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21381_ VGND VPWR _01426_ _06150_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_31_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20332_ VGND VPWR _00935_ _05592_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_259_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23120_ VPWR VGND VGND VPWR _07039_ _03488_ _03490_ sky130_fd_sc_hd__nand2_2
XFILLER_0_226_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23051_ VGND VPWR VGND VPWR _03254_ _03795_ _03255_ _03257_ _06998_ _06892_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_12_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20263_ VGND VPWR VPWR VGND _05546_ _02410_ keymem.key_mem\[9\]\[19\] _05556_ sky130_fd_sc_hd__mux2_2
XFILLER_0_101_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1061 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22002_ VGND VPWR VGND VPWR _06481_ keymem.key_mem_we _03194_ _06475_ _01716_ sky130_fd_sc_hd__a31o_2
X_20194_ VGND VPWR VPWR VGND _05515_ _03592_ keymem.key_mem\[10\]\[116\] _05518_ sky130_fd_sc_hd__mux2_2
XFILLER_0_122_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23953_ VGND VPWR VPWR VGND clk _00446_ reset_n keymem.key_mem\[13\]\[74\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_97_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_192_1227 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_157_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22904_ VGND VPWR VGND VPWR _06908_ _11108_ _03860_ _06884_ _11147_ sky130_fd_sc_hd__a211o_2
XFILLER_0_223_260 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23884_ VGND VPWR VPWR VGND clk _00377_ reset_n keymem.key_mem\[13\]\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_196_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_93_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25623_ VGND VPWR VPWR VGND clk _02116_ reset_n keymem.key_mem\[0\]\[80\] sky130_fd_sc_hd__dfrtp_2
X_22835_ VPWR VGND VPWR VGND _06866_ keymem.rcon_reg\[0\] keymem.rcon_logic.tmp_rcon\[0\]
+ sky130_fd_sc_hd__or2_2
XFILLER_0_168_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25554_ VGND VPWR VPWR VGND clk _02047_ reset_n keymem.key_mem\[0\]\[11\] sky130_fd_sc_hd__dfrtp_2
X_22766_ VGND VPWR VPWR VGND _06833_ keymem.key_mem\[0\]\[80\] _03330_ _06846_ sky130_fd_sc_hd__mux2_2
X_24505_ VGND VPWR VPWR VGND clk _00998_ reset_n keymem.key_mem\[9\]\[114\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21717_ VGND VPWR VPWR VGND _06319_ _03161_ keymem.key_mem\[4\]\[61\] _06328_ sky130_fd_sc_hd__mux2_2
X_25485_ VGND VPWR VPWR VGND clk _01978_ reset_n keymem.key_mem\[1\]\[70\] sky130_fd_sc_hd__dfrtp_2
X_22697_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[38\] _06790_ _06789_ _04931_ _02074_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_240_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_107_1_Right_708 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12450_ VPWR VGND VPWR VGND keymem.key_mem\[8\]\[30\] _07752_ keymem.key_mem\[1\]\[30\]
+ _07557_ _08023_ sky130_fd_sc_hd__a22o_2
X_24436_ VGND VPWR VPWR VGND clk _00929_ reset_n keymem.key_mem\[9\]\[45\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_168_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_111_2_Right_183 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21648_ VGND VPWR VPWR VGND _06286_ _02786_ keymem.key_mem\[4\]\[28\] _06292_ sky130_fd_sc_hd__mux2_2
XFILLER_0_30_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_243 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_168_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12381_ VGND VPWR VGND VPWR _07960_ _07958_ keymem.key_mem\[8\]\[24\] _07959_ _07572_
+ sky130_fd_sc_hd__a211o_2
X_24367_ VGND VPWR VPWR VGND clk _00860_ reset_n keymem.key_mem\[10\]\[104\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_34_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21579_ VGND VPWR VPWR VGND _06116_ _03654_ keymem.key_mem\[5\]\[125\] _06254_ sky130_fd_sc_hd__mux2_2
XFILLER_0_50_725 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14120_ VPWR VGND VGND VPWR _09422_ _09591_ _09354_ sky130_fd_sc_hd__nor2_2
X_23318_ VPWR VGND VGND VPWR _07198_ _07194_ _07196_ sky130_fd_sc_hd__nand2_2
XFILLER_0_65_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24298_ VGND VPWR VPWR VGND clk _00791_ reset_n keymem.key_mem\[10\]\[35\] sky130_fd_sc_hd__dfrtp_2
X_14051_ VGND VPWR _09523_ _09510_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23249_ VPWR VGND VPWR VGND _07135_ block[4] _03957_ enc_block.block_w2_reg\[4\]
+ _03952_ _07136_ sky130_fd_sc_hd__a221o_2
XFILLER_0_104_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_1161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_247_831 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13002_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[83\] _08449_ _08521_ _08517_ _08522_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_24_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_105_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_219_555 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_140_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17810_ VPWR VGND VPWR VGND _03170_ _03802_ keymem.prev_key0_reg\[62\] _03788_ _00203_
+ sky130_fd_sc_hd__a22o_2
X_18790_ _04640_ _04642_ _03982_ _04641_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_101_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17741_ VGND VPWR VPWR VGND _03723_ _02915_ keymem.prev_key0_reg\[37\] _03759_ sky130_fd_sc_hd__mux2_2
X_14953_ VGND VPWR VGND VPWR enc_block.block_w2_reg\[12\] _09269_ _09021_ _10415_
+ _10417_ _10416_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_101_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_175_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13904_ VGND VPWR VPWR VGND _09363_ _09375_ _09373_ _09376_ sky130_fd_sc_hd__or3_2
XFILLER_0_76_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17672_ VGND VPWR VPWR VGND _03691_ key[144] keymem.prev_key1_reg\[16\] _03711_ sky130_fd_sc_hd__mux2_2
X_14884_ VGND VPWR VPWR VGND _10026_ _10348_ _10022_ _10349_ sky130_fd_sc_hd__or3_2
XFILLER_0_72_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_255_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19411_ VGND VPWR VGND VPWR _05101_ keymem.key_mem_we _10194_ _05093_ _00505_ sky130_fd_sc_hd__a31o_2
X_16623_ VGND VPWR VGND VPWR _02777_ _02776_ _02778_ _02779_ sky130_fd_sc_hd__a21o_2
X_13835_ VGND VPWR VGND VPWR _09307_ _09279_ _09278_ keymem.prev_key1_reg\[30\] _08989_
+ _08983_ sky130_fd_sc_hd__a32o_2
XFILLER_0_159_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_202_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19342_ VGND VPWR _00482_ _05055_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16554_ VGND VPWR VGND VPWR _02710_ _02711_ _02713_ _02709_ sky130_fd_sc_hd__nand3_2
XFILLER_0_43_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_184 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13766_ VGND VPWR VGND VPWR _09193_ _09237_ _09238_ _09183_ _09214_ sky130_fd_sc_hd__nor4_2
XFILLER_0_202_499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15505_ VGND VPWR _09512_ key[12] _10965_ _08936_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_112_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12717_ VGND VPWR _08265_ _07540_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19273_ VGND VPWR VPWR VGND _04993_ _05010_ keymem.key_mem\[13\]\[86\] _05011_ sky130_fd_sc_hd__mux2_2
X_16485_ _02643_ _02646_ keymem.prev_key0_reg\[23\] _02644_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_151_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13697_ VGND VPWR VGND VPWR _09146_ _09095_ _09167_ _09169_ sky130_fd_sc_hd__a21o_2
X_18224_ VPWR VGND VPWR VGND _04131_ block[110] _03980_ enc_block.block_w2_reg\[14\]
+ _03978_ _04132_ sky130_fd_sc_hd__a221o_2
XFILLER_0_112_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15436_ VPWR VGND _10897_ _10896_ keymem.prev_key0_reg\[11\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_5_605 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12648_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[49\] _07695_ keymem.key_mem\[4\]\[49\]
+ _07693_ _08202_ sky130_fd_sc_hd__a22o_2
XFILLER_0_186_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18155_ VPWR VGND VPWR VGND _04069_ _03983_ _04067_ sky130_fd_sc_hd__or2_2
XFILLER_0_147_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_182_395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15367_ VGND VPWR _10829_ keymem.prev_key1_reg\[74\] _10828_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12579_ VPWR VGND VPWR VGND _08139_ keymem.key_mem\[10\]\[42\] _07785_ keymem.key_mem\[8\]\[42\]
+ _07655_ _08140_ sky130_fd_sc_hd__a221o_2
XFILLER_0_83_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_104_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17106_ VPWR VGND _03222_ _03221_ keymem.prev_key0_reg\[68\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_4_159 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14318_ VGND VPWR VGND VPWR _09618_ _09361_ _09781_ _09783_ _09788_ _09787_ sky130_fd_sc_hd__a2111o_2
X_18086_ VPWR VGND VGND VPWR _04005_ _04006_ _03993_ sky130_fd_sc_hd__nor2_2
XFILLER_0_262_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15298_ VGND VPWR VGND VPWR _10668_ _10667_ _10760_ _10498_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_83_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17037_ VPWR VGND VPWR VGND _03160_ _10086_ _03157_ _03158_ _03159_ _10096_ sky130_fd_sc_hd__o311a_2
X_14249_ VPWR VGND VPWR VGND _09720_ key[1] _09719_ sky130_fd_sc_hd__or2_2
XFILLER_0_262_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_493 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_123_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_352 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_225_514 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18988_ VPWR VGND _04820_ _04819_ enc_block.round_key\[56\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_193_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17939_ VGND VPWR _00244_ _03890_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_20_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20950_ VGND VPWR VPWR VGND _05912_ _05006_ keymem.key_mem\[7\]\[84\] _05922_ sky130_fd_sc_hd__mux2_2
XFILLER_0_234_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_205_271 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19609_ VGND VPWR _00597_ _05207_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_5_Right_5 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20881_ VGND VPWR VPWR VGND _05880_ _04958_ keymem.key_mem\[7\]\[52\] _05885_ sky130_fd_sc_hd__mux2_2
XFILLER_0_36_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_7_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22620_ VGND VPWR VPWR VGND _06779_ keymem.key_mem\[0\]\[0\] _09537_ _06780_ sky130_fd_sc_hd__mux2_2
XFILLER_0_152_1266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22551_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[77\] _06754_ _06753_ _04995_ _01985_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_8_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_90_102 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_130_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21502_ VGND VPWR VPWR VGND _06209_ _03401_ keymem.key_mem\[5\]\[88\] _06214_ sky130_fd_sc_hd__mux2_2
XFILLER_0_8_454 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25270_ VGND VPWR VPWR VGND clk _01763_ reset_n keymem.key_mem\[3\]\[111\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_210 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_63_349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22482_ VGND VPWR _01943_ _06734_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_118_278 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24221_ VGND VPWR VPWR VGND clk _00714_ reset_n keymem.key_mem\[11\]\[86\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_267_1397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21433_ VGND VPWR VPWR VGND _06173_ _03099_ keymem.key_mem\[5\]\[55\] _06178_ sky130_fd_sc_hd__mux2_2
XFILLER_0_12_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21364_ VGND VPWR VPWR VGND _06140_ _02607_ keymem.key_mem\[5\]\[22\] _06142_ sky130_fd_sc_hd__mux2_2
X_24152_ VGND VPWR VPWR VGND clk _00645_ reset_n keymem.key_mem\[11\]\[17\] sky130_fd_sc_hd__dfrtp_2
X_20315_ VGND VPWR _00927_ _05583_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23103_ VGND VPWR VPWR VGND _06992_ _07028_ keymem.prev_key1_reg\[93\] _07029_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_241_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24083_ VGND VPWR VPWR VGND clk _00576_ reset_n keymem.key_mem\[12\]\[76\] sky130_fd_sc_hd__dfrtp_2
X_21295_ VGND VPWR VPWR VGND _06098_ _03613_ keymem.key_mem\[6\]\[119\] _06104_ sky130_fd_sc_hd__mux2_2
XFILLER_0_141_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_248_639 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_1481 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_229_831 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23034_ VGND VPWR VGND VPWR _02243_ _06986_ _06954_ keymem.prev_key1_reg\[66\] sky130_fd_sc_hd__o21a_2
X_20246_ VGND VPWR _00894_ _05547_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20177_ VGND VPWR VPWR VGND _05504_ _03543_ keymem.key_mem\[10\]\[108\] _05509_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_186_1_Left_453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_243_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_154_2_Left_625 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24985_ VGND VPWR VPWR VGND clk _01478_ reset_n keymem.key_mem\[5\]\[82\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_243_355 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_235_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23936_ VGND VPWR VPWR VGND clk _00429_ reset_n keymem.key_mem\[13\]\[57\] sky130_fd_sc_hd__dfrtp_2
X_11950_ VPWR VGND VPWR VGND keymem.key_mem\[4\]\[0\] _07552_ keymem.key_mem\[2\]\[0\]
+ _07547_ _07553_ sky130_fd_sc_hd__a22o_2
XFILLER_0_197_922 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_157_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11881_ VGND VPWR result[107] _07504_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23867_ VGND VPWR VPWR VGND clk _00360_ reset_n enc_block.block_w2_reg\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13620_ VGND VPWR VGND VPWR _09090_ _09091_ _09036_ _09087_ _09085_ _09092_ sky130_fd_sc_hd__o32a_2
X_25606_ VGND VPWR VPWR VGND clk _02099_ reset_n keymem.key_mem\[0\]\[63\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_233_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22818_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[117\] _06860_ _06859_ _05069_ _02153_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_168_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23798_ VGND VPWR VPWR VGND clk _00291_ reset_n enc_block.block_w0_reg\[17\] sky130_fd_sc_hd__dfrtp_2
X_13551_ enc_block.sword_ctr_reg\[1\] _09023_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[0\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_109_212 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25537_ VGND VPWR VPWR VGND clk _02030_ reset_n keymem.key_mem\[1\]\[122\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22749_ VGND VPWR _06840_ _03227_ _02104_ _06839_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_66_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_251_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_327 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12502_ VGND VPWR VGND VPWR _07691_ keymem.key_mem\[3\]\[35\] _08066_ _08068_ _08070_
+ _08069_ sky130_fd_sc_hd__a2111o_2
X_16270_ VPWR VGND VPWR VGND _02432_ _02433_ _02434_ _02385_ _02431_ sky130_fd_sc_hd__or4b_2
XFILLER_0_66_187 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13482_ VGND VPWR _08954_ _08938_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25468_ VGND VPWR VPWR VGND clk _01961_ reset_n keymem.key_mem\[1\]\[53\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_246_1415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15221_ VGND VPWR VGND VPWR _10480_ _10574_ _10608_ _10612_ _10684_ sky130_fd_sc_hd__o22a_2
XPHY_EDGE_ROW_108_1_Right_709 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24419_ VGND VPWR VPWR VGND clk _00912_ reset_n keymem.key_mem\[9\]\[28\] sky130_fd_sc_hd__dfrtp_2
X_12433_ VGND VPWR VGND VPWR _07800_ keymem.key_mem\[1\]\[29\] _08004_ _08006_ _08007_
+ _07663_ sky130_fd_sc_hd__a2111o_2
XPHY_EDGE_ROW_112_2_Right_184 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_120_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25399_ VGND VPWR VPWR VGND clk _01892_ reset_n keymem.key_mem\[2\]\[112\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_585 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15152_ VGND VPWR VGND VPWR _10616_ _10615_ _10614_ _10613_ _10607_ sky130_fd_sc_hd__and4_2
XFILLER_0_50_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12364_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[23\] _07596_ keymem.key_mem\[4\]\[23\]
+ _07551_ _07944_ sky130_fd_sc_hd__a22o_2
XFILLER_0_209_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14103_ _09370_ _09574_ _09247_ _09573_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_65_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15083_ VGND VPWR _10547_ _10546_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_26_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19960_ VGND VPWR VPWR VGND _05389_ _10194_ keymem.key_mem\[10\]\[5\] _05395_ sky130_fd_sc_hd__mux2_2
X_12295_ VPWR VGND VPWR VGND _07880_ keymem.key_mem\[6\]\[17\] _07818_ keymem.key_mem\[2\]\[17\]
+ _07733_ _07881_ sky130_fd_sc_hd__a221o_2
XFILLER_0_267_959 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18911_ VPWR VGND _04751_ _04750_ enc_block.round_key\[48\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_14034_ _09429_ _09506_ _09240_ _09505_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_201_1009 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_238_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_129_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19891_ VGND VPWR VPWR VGND _05350_ keymem.key_mem\[11\]\[102\] _03506_ _05357_ sky130_fd_sc_hd__mux2_2
X_18842_ VPWR VGND VGND VPWR _04688_ _04689_ enc_block.round_key\[41\] sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_86_2_Left_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18773_ VPWR VGND _04626_ enc_block.block_w2_reg\[27\] enc_block.block_w3_reg\[19\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_15985_ VGND VPWR _11441_ keymem.prev_key0_reg\[112\] _11440_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_234_344 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_179_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_145_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_250_826 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14936_ VGND VPWR VGND VPWR enc_block.block_w1_reg\[10\] _08947_ _09021_ _10398_
+ _10400_ _10399_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_261_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_234_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17724_ VGND VPWR VGND VPWR _03732_ keymem.prev_key1_reg\[30\] _03749_ _03733_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_89_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14867_ VPWR VGND VPWR VGND _10331_ _10019_ _09803_ _09189_ _09012_ _10332_ sky130_fd_sc_hd__a221o_2
XFILLER_0_72_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17655_ VGND VPWR _00151_ _03699_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_37_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13818_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[28\] _08989_ _09290_ _08983_ _09288_
+ _09289_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_225_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16606_ VPWR VGND VPWR VGND _02763_ _10325_ _02760_ _02761_ _02762_ _10281_ sky130_fd_sc_hd__o311a_2
XFILLER_0_212_1127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17586_ _03644_ _03646_ _09533_ _03645_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_14798_ VGND VPWR keymem.prev_key0_reg\[102\] _10230_ _10264_ _10262_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_212_1138 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19325_ VGND VPWR VPWR VGND _05025_ _05043_ keymem.key_mem\[13\]\[105\] _05044_ sky130_fd_sc_hd__mux2_2
X_16537_ VPWR VGND VGND VPWR keymem.prev_key0_reg\[121\] _02695_ _07387_ _02693_ _02694_
+ _02696_ sky130_fd_sc_hd__a311o_2
X_13749_ VGND VPWR _09221_ _09200_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_35_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16468_ VGND VPWR VGND VPWR _11218_ _11330_ _11235_ _11403_ _02629_ sky130_fd_sc_hd__o22a_2
X_19256_ VGND VPWR VGND VPWR _05000_ keymem.key_mem_we _03322_ _04999_ _00451_ sky130_fd_sc_hd__a31o_2
XFILLER_0_112_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15419_ VPWR VGND VGND VPWR _10668_ _10511_ _10609_ _10455_ _10880_ _10549_ sky130_fd_sc_hd__o221a_2
X_18207_ VPWR VGND VGND VPWR _04116_ _04117_ _04041_ sky130_fd_sc_hd__nor2_2
XFILLER_0_182_170 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_72_168 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19187_ VGND VPWR VPWR VGND _04951_ _04958_ keymem.key_mem\[13\]\[52\] _04959_ sky130_fd_sc_hd__mux2_2
X_16399_ VPWR VGND VGND VPWR _02424_ _02524_ _02560_ _02561_ sky130_fd_sc_hd__nor3_2
XFILLER_0_147_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_371 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_14_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18138_ VPWR VGND VPWR VGND _04053_ _04040_ _04051_ enc_block.block_w0_reg\[6\] _03976_
+ _00280_ sky130_fd_sc_hd__a221o_2
XFILLER_0_83_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_53_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18069_ VPWR VGND VPWR VGND _03989_ block[97] _03980_ enc_block.block_w3_reg\[1\]
+ _03978_ _03990_ sky130_fd_sc_hd__a221o_2
XFILLER_0_123_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_44_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_292 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20100_ VGND VPWR _00827_ _05468_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21080_ VGND VPWR _01284_ _05991_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_95_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20031_ VGND VPWR _00794_ _05432_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_186_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_158_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_256_1043 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_119_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_225_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24770_ VGND VPWR VPWR VGND clk _01263_ reset_n keymem.key_mem\[7\]\[123\] sky130_fd_sc_hd__dfrtp_2
X_21982_ VGND VPWR VPWR VGND _06462_ _04963_ keymem.key_mem\[3\]\[55\] _06471_ sky130_fd_sc_hd__mux2_2
XFILLER_0_94_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23721_ keymem.prev_key0_reg\[77\] clk _00218_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20933_ VGND VPWR VPWR VGND _05912_ _04992_ keymem.key_mem\[7\]\[76\] _05913_ sky130_fd_sc_hd__mux2_2
XFILLER_0_7_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_16_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23652_ keymem.prev_key0_reg\[8\] clk _00149_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_7_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20864_ VGND VPWR VPWR VGND _05867_ _04943_ keymem.key_mem\[7\]\[44\] _05876_ sky130_fd_sc_hd__mux2_2
XFILLER_0_165_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22603_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[113\] _06777_ _06776_ _05060_ _02021_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_7_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23583_ VGND VPWR VPWR VGND clk _00084_ reset_n keymem.key_mem\[14\]\[72\] sky130_fd_sc_hd__dfrtp_2
X_20795_ VPWR VGND keymem.key_mem\[7\]\[12\] _05839_ _05830_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_63_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_63_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25322_ VGND VPWR VPWR VGND clk _01815_ reset_n keymem.key_mem\[2\]\[35\] sky130_fd_sc_hd__dfrtp_2
X_22534_ VGND VPWR VPWR VGND _06750_ keymem.key_mem\[1\]\[67\] _03217_ _06755_ sky130_fd_sc_hd__mux2_2
XFILLER_0_187_1159 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_64_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_267_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1003 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_169_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25253_ VGND VPWR VPWR VGND clk _01746_ reset_n keymem.key_mem\[3\]\[94\] sky130_fd_sc_hd__dfrtp_2
X_22465_ VGND VPWR VPWR VGND _06726_ keymem.key_mem\[1\]\[26\] _02743_ _06727_ sky130_fd_sc_hd__mux2_2
XFILLER_0_165_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_585 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24204_ VGND VPWR VPWR VGND clk _00697_ reset_n keymem.key_mem\[11\]\[69\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_66_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21416_ VGND VPWR VPWR VGND _06162_ _03024_ keymem.key_mem\[5\]\[47\] _06169_ sky130_fd_sc_hd__mux2_2
XFILLER_0_60_842 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_126_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25184_ VGND VPWR VPWR VGND clk _01677_ reset_n keymem.key_mem\[3\]\[25\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_228_1189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22396_ VGND VPWR _01902_ _06689_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_165_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24135_ VGND VPWR VPWR VGND clk _00628_ reset_n keymem.key_mem\[11\]\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_886 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21347_ VGND VPWR VPWR VGND _06128_ _11098_ keymem.key_mem\[5\]\[14\] _06133_ sky130_fd_sc_hd__mux2_2
XFILLER_0_27_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_292 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_206_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24066_ VGND VPWR VPWR VGND clk _00559_ reset_n keymem.key_mem\[12\]\[59\] sky130_fd_sc_hd__dfrtp_2
X_12080_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[4\] _07591_ keymem.key_mem\[4\]\[4\]
+ _07550_ _07679_ sky130_fd_sc_hd__a22o_2
X_21278_ VGND VPWR VPWR VGND _06087_ _03560_ keymem.key_mem\[6\]\[111\] _06095_ sky130_fd_sc_hd__mux2_2
X_23017_ VGND VPWR VPWR VGND _02235_ _03123_ _03128_ _06925_ _06977_ sky130_fd_sc_hd__o31a_2
XFILLER_0_217_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20229_ VGND VPWR _00886_ _05538_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_102_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15770_ VGND VPWR _11226_ _11225_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_176_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12982_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[81\] _08449_ _08503_ _08499_ _08504_
+ sky130_fd_sc_hd__o22a_2
X_24968_ VGND VPWR VPWR VGND clk _01461_ reset_n keymem.key_mem\[5\]\[65\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_73_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14721_ VGND VPWR VPWR VGND _10147_ _10187_ _09932_ _10188_ sky130_fd_sc_hd__or3_2
XFILLER_0_137_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23919_ VGND VPWR VPWR VGND clk _00412_ reset_n keymem.key_mem\[13\]\[40\] sky130_fd_sc_hd__dfrtp_2
X_11933_ VGND VPWR _07536_ _07535_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_19_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_73_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24899_ VGND VPWR VPWR VGND clk _01392_ reset_n keymem.key_mem\[6\]\[124\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_34_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17440_ VGND VPWR _00116_ _03519_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_213_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14652_ VPWR VGND VPWR VGND _09915_ _10118_ _10119_ _09595_ _09760_ sky130_fd_sc_hd__or4b_2
XFILLER_0_19_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11864_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[3\] dec_new_block\[99\]
+ _07496_ sky130_fd_sc_hd__mux2_2
XFILLER_0_39_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_170_1163 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_196_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13603_ VPWR VGND VGND VPWR _09038_ _09055_ _09074_ _09075_ sky130_fd_sc_hd__nor3_2
XFILLER_0_213_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17371_ VGND VPWR _03460_ _03459_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14583_ VPWR VGND VPWR VGND _09465_ _09596_ _10051_ _10049_ _10050_ sky130_fd_sc_hd__or4b_2
XFILLER_0_39_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11795_ VGND VPWR result[64] _07461_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_131_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16322_ VPWR VGND VPWR VGND _02485_ keymem.prev_key1_reg\[117\] sky130_fd_sc_hd__inv_2
X_19110_ VGND VPWR VGND VPWR _04910_ keymem.key_mem_we _02661_ _04908_ _00395_ sky130_fd_sc_hd__a31o_2
X_13534_ VPWR VGND VPWR VGND _08982_ _09005_ _08991_ _09001_ _09006_ sky130_fd_sc_hd__or4_2
XFILLER_0_40_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_198 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19041_ VPWR VGND VGND VPWR _04600_ _04867_ _04292_ sky130_fd_sc_hd__nor2_2
X_16253_ VPWR VGND VPWR VGND _11611_ _02416_ _02413_ _11566_ _02417_ sky130_fd_sc_hd__or4_2
XFILLER_0_36_861 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_246_1223 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13465_ VGND VPWR _08937_ _08936_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_10_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15204_ VGND VPWR _10667_ _10437_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_35_382 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12416_ VGND VPWR VGND VPWR _07992_ _07619_ keymem.key_mem\[3\]\[27\] _07989_ _07991_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_152_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16184_ VPWR VGND VGND VPWR _11425_ _02348_ _02349_ sky130_fd_sc_hd__or2b_2
XFILLER_0_35_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_113_2_Right_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_853 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13396_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[123\] _07596_ keymem.key_mem\[13\]\[123\]
+ _07587_ _08876_ sky130_fd_sc_hd__a22o_2
XFILLER_0_144_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15135_ VGND VPWR VGND VPWR _10528_ _10527_ _10599_ _10508_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_80_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_105_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12347_ VGND VPWR _07929_ _07539_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_10_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_267_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15066_ VGND VPWR _10530_ _10529_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19943_ VGND VPWR VPWR VGND _05246_ keymem.key_mem\[11\]\[127\] _03668_ _05384_ sky130_fd_sc_hd__mux2_2
XFILLER_0_10_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_220_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12278_ VGND VPWR _07865_ _07560_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_267_778 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_254_406 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14017_ VPWR VGND VGND VPWR _09489_ _09361_ _09362_ sky130_fd_sc_hd__nand2_2
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19874_ VGND VPWR VPWR VGND _05339_ keymem.key_mem\[11\]\[94\] _03452_ _05348_ sky130_fd_sc_hd__mux2_2
X_18825_ VPWR VGND VGND VPWR _04654_ _04674_ _04062_ sky130_fd_sc_hd__nor2_2
XFILLER_0_120_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18756_ VPWR VGND VPWR VGND _04610_ block[33] _04576_ enc_block.block_w1_reg\[1\]
+ _04543_ _04611_ sky130_fd_sc_hd__a221o_2
X_15968_ VPWR VGND VPWR VGND _11421_ _11423_ _11424_ _11416_ _11418_ sky130_fd_sc_hd__or4b_2
XFILLER_0_250_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_222_336 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17707_ VGND VPWR _03737_ _02647_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_76_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14919_ VPWR VGND VGND VPWR _10383_ key[136] _09544_ sky130_fd_sc_hd__nand2_2
X_15899_ VPWR VGND VGND VPWR _11325_ _11355_ _11210_ sky130_fd_sc_hd__nor2_2
X_18687_ VPWR VGND _04549_ _04548_ enc_block.round_key\[90\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_8_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_231_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17638_ VGND VPWR VPWR VGND _03681_ _03687_ keymem.prev_key0_reg\[5\] _03688_ sky130_fd_sc_hd__mux2_2
XFILLER_0_59_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1093 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_187_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_147_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_231_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17569_ VPWR VGND VPWR VGND _03631_ key[250] _09927_ sky130_fd_sc_hd__or2_2
XFILLER_0_18_327 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19308_ VGND VPWR _00471_ _05032_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_85_293 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20580_ VGND VPWR VPWR VGND _05714_ _02964_ keymem.key_mem\[8\]\[41\] _05723_ sky130_fd_sc_hd__mux2_2
XFILLER_0_45_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_45_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_61_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19239_ VGND VPWR VGND VPWR _03277_ _03276_ _04989_ _08921_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_45_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_243 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_382 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_42_842 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22250_ VGND VPWR _01832_ _06613_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21201_ VPWR VGND VGND VPWR _06055_ keymem.key_mem\[6\]\[74\] _05985_ sky130_fd_sc_hd__nand2_2
XFILLER_0_147_1187 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_48_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22181_ VGND VPWR VPWR VGND _06565_ _02479_ keymem.key_mem\[2\]\[20\] _06577_ sky130_fd_sc_hd__mux2_2
XFILLER_0_2_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1042 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21132_ VGND VPWR VPWR VGND _06018_ _02964_ keymem.key_mem\[6\]\[41\] _06019_ sky130_fd_sc_hd__mux2_2
XFILLER_0_1_460 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_111_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21063_ VGND VPWR VPWR VGND _05972_ _10746_ keymem.key_mem\[6\]\[9\] _05982_ sky130_fd_sc_hd__mux2_2
XFILLER_0_160_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20014_ VGND VPWR _00786_ _05423_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24822_ VGND VPWR VPWR VGND clk _01315_ reset_n keymem.key_mem\[6\]\[47\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24753_ VGND VPWR VPWR VGND clk _01246_ reset_n keymem.key_mem\[7\]\[106\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21965_ VGND VPWR VGND VPWR _06461_ keymem.key_mem_we _03025_ _06446_ _01699_ sky130_fd_sc_hd__a31o_2
X_23704_ keymem.prev_key0_reg\[60\] clk _00201_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20916_ VPWR VGND VGND VPWR _05904_ keymem.key_mem\[7\]\[68\] _05824_ sky130_fd_sc_hd__nand2_2
XFILLER_0_90_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24684_ VGND VPWR VPWR VGND clk _01177_ reset_n keymem.key_mem\[7\]\[37\] sky130_fd_sc_hd__dfrtp_2
X_21896_ VGND VPWR VGND VPWR _06424_ keymem.key_mem_we _11149_ _06420_ _01667_ sky130_fd_sc_hd__a31o_2
X_23635_ VGND VPWR VPWR VGND clk _00136_ reset_n keymem.key_mem\[14\]\[124\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_193_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20847_ VGND VPWR _05867_ _05819_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_162_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23566_ VGND VPWR VPWR VGND clk _00067_ reset_n keymem.key_mem\[14\]\[55\] sky130_fd_sc_hd__dfrtp_2
X_20778_ VGND VPWR VGND VPWR _05829_ keymem.key_mem_we _10099_ _05821_ _01144_ sky130_fd_sc_hd__a31o_2
X_25305_ VGND VPWR VPWR VGND clk _01798_ reset_n keymem.key_mem\[2\]\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_64_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22517_ VGND VPWR VPWR VGND _06739_ keymem.key_mem\[1\]\[59\] _03140_ _06746_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_360 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23497_ VGND VPWR _07357_ enc_block.block_w0_reg\[23\] _07148_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_134_343 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_165_1232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_140 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_134_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25236_ VGND VPWR VPWR VGND clk _01729_ reset_n keymem.key_mem\[3\]\[77\] sky130_fd_sc_hd__dfrtp_2
X_13250_ VPWR VGND VPWR VGND _08744_ keymem.key_mem\[10\]\[108\] _07909_ keymem.key_mem\[1\]\[108\]
+ _07715_ _08745_ sky130_fd_sc_hd__a221o_2
XFILLER_0_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_1059 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22448_ VGND VPWR VPWR VGND _06715_ keymem.key_mem\[1\]\[18\] _02340_ _06718_ sky130_fd_sc_hd__mux2_2
XFILLER_0_126_1216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_66_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12201_ VGND VPWR VGND VPWR _07793_ keymem.key_mem\[0\]\[10\] _07792_ _07784_ _07777_
+ _07794_ sky130_fd_sc_hd__o32a_2
X_13181_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[101\] _07724_ keymem.key_mem\[7\]\[101\]
+ _07702_ _08683_ sky130_fd_sc_hd__a22o_2
X_25167_ VGND VPWR VPWR VGND clk _01660_ reset_n keymem.key_mem\[3\]\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22379_ VGND VPWR VPWR VGND _06680_ _03580_ keymem.key_mem\[2\]\[114\] _06681_ sky130_fd_sc_hd__mux2_2
XFILLER_0_66_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24118_ VGND VPWR VPWR VGND clk _00611_ reset_n keymem.key_mem\[12\]\[111\] sky130_fd_sc_hd__dfrtp_2
X_12132_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[6\] _07645_ _07728_ _07720_ _07729_
+ sky130_fd_sc_hd__o22a_2
X_25098_ VGND VPWR VPWR VGND clk _01591_ reset_n keymem.key_mem\[4\]\[67\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_102_284 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16940_ VGND VPWR VPWR VGND _10091_ key[180] keymem.prev_key1_reg\[52\] _03072_ sky130_fd_sc_hd__mux2_2
X_12063_ VGND VPWR _07663_ _07662_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24049_ VGND VPWR VPWR VGND clk _00542_ reset_n keymem.key_mem\[12\]\[42\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_257_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1074 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16871_ VGND VPWR _02866_ key[46] _03009_ _10189_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_99_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18610_ VGND VPWR _04480_ enc_block.block_w0_reg\[2\] _04479_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15822_ VPWR VGND VGND VPWR _11278_ _11263_ _11174_ sky130_fd_sc_hd__nand2_2
X_19590_ VGND VPWR _00588_ _05197_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_35_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1082 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_137_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_149_1_Left_416 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15753_ VPWR VGND VPWR VGND _11206_ _11208_ _11207_ _11187_ _11209_ sky130_fd_sc_hd__or4_2
X_18541_ VPWR VGND VPWR VGND _04418_ _04343_ _04417_ sky130_fd_sc_hd__or2_2
XFILLER_0_73_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12965_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[80\] _07599_ keymem.key_mem\[10\]\[80\]
+ _07560_ _08488_ sky130_fd_sc_hd__a22o_2
XFILLER_0_99_374 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_137_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11916_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[29\] dec_new_block\[125\]
+ _07522_ sky130_fd_sc_hd__mux2_2
X_14704_ VGND VPWR VGND VPWR _09079_ _09126_ _09121_ _09115_ _10171_ sky130_fd_sc_hd__o22a_2
X_15684_ VPWR VGND VGND VPWR _11120_ _11135_ _11138_ _11140_ _11141_ sky130_fd_sc_hd__and4b_2
XFILLER_0_34_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18472_ VPWR VGND _04356_ _04355_ _04354_ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_231_188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_38_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12896_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[73\] _07702_ keymem.key_mem\[6\]\[73\]
+ _07656_ _08426_ sky130_fd_sc_hd__a22o_2
XFILLER_0_213_1233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17423_ VPWR VGND _09533_ _03505_ _03504_ VPWR VGND sky130_fd_sc_hd__and2_2
X_14635_ VPWR VGND VPWR VGND _10102_ _10101_ sky130_fd_sc_hd__inv_2
X_11847_ VGND VPWR result[90] _07487_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_129_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_265 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14566_ _09478_ _10034_ _09550_ _09364_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_67_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17354_ VGND VPWR VPWR VGND _03384_ keymem.key_mem\[14\]\[93\] _03444_ _03445_ sky130_fd_sc_hd__mux2_2
X_11778_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[24\] dec_new_block\[56\]
+ _07453_ sky130_fd_sc_hd__mux2_2
XFILLER_0_51_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13517_ VGND VPWR _08989_ _08954_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16305_ VPWR VGND _02469_ keymem.prev_key1_reg\[52\] keymem.prev_key1_reg\[20\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
X_17285_ VPWR VGND VPWR VGND _03382_ _03379_ _03378_ key[214] _03366_ _03383_ sky130_fd_sc_hd__a221o_2
XFILLER_0_15_319 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14497_ VPWR VGND VPWR VGND _09956_ _09965_ _09960_ _09055_ _09966_ sky130_fd_sc_hd__or4_2
X_19024_ VPWR VGND _04852_ _04851_ enc_block.round_key\[60\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_109_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16236_ VGND VPWR VPWR VGND _02400_ _02398_ _02397_ _02401_ sky130_fd_sc_hd__mux2_2
X_13448_ VPWR VGND VGND VPWR _07389_ _00003_ _08922_ sky130_fd_sc_hd__nor2_2
XFILLER_0_148_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_84_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_352 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16167_ VGND VPWR VGND VPWR _11619_ keymem.round_ctr_reg\[0\] _11620_ _11621_ sky130_fd_sc_hd__a21o_2
XPHY_EDGE_ROW_114_2_Right_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_374 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13379_ VGND VPWR VGND VPWR _07778_ keymem.key_mem\[3\]\[121\] _08858_ _08860_ _08861_
+ _08736_ sky130_fd_sc_hd__a2111o_2
X_15118_ VPWR VGND VPWR VGND _10571_ _10581_ _10577_ _10561_ _10582_ sky130_fd_sc_hd__or4_2
XFILLER_0_45_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16098_ VPWR VGND VPWR VGND _11552_ _11551_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15049_ VGND VPWR _10513_ _10503_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_259_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19926_ VGND VPWR _00746_ _05375_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_167_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19857_ VGND VPWR _05339_ _05242_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_254_269 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_208_664 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18808_ VGND VPWR _04658_ enc_block.block_w1_reg\[5\] _04657_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_257_1160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_208_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19788_ VGND VPWR _05303_ _05246_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_155_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18739_ VPWR VGND VPWR VGND _04595_ _04591_ _04593_ sky130_fd_sc_hd__or2_2
XFILLER_0_116_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21750_ VGND VPWR _01600_ _06345_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_750 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_116_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20701_ VGND VPWR _01110_ _05786_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_8_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21681_ VGND VPWR _01567_ _06309_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_175_232 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_70_1_Left_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_231_1377 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_945 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23420_ VGND VPWR VGND VPWR _07289_ _04149_ _07095_ _07290_ enc_block.block_w3_reg\[21\]
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_50_1152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20632_ VGND VPWR _01077_ _05750_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_266_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_606 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23351_ VPWR VGND VGND VPWR _07228_ enc_block.round_key\[14\] _07227_ sky130_fd_sc_hd__nand2_2
XFILLER_0_116_321 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_195_1_Left_462 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_128_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20563_ VGND VPWR _05714_ _05679_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_11_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_91 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22302_ VGND VPWR _01857_ _06640_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_163_2_Left_634 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_116_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_127_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23282_ VPWR VGND VPWR VGND _07165_ _04874_ _07164_ enc_block.block_w3_reg\[7\] _07115_
+ _02312_ sky130_fd_sc_hd__a221o_2
XFILLER_0_166_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20494_ VGND VPWR _01012_ _05677_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_127_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25021_ VGND VPWR VPWR VGND clk _01514_ reset_n keymem.key_mem\[5\]\[118\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22233_ VGND VPWR _01824_ _06604_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_225_1159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_160_1_Right_761 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22164_ VGND VPWR _06568_ _10913_ _01791_ _06567_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_258_564 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_219_918 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21115_ VGND VPWR VPWR VGND _06007_ _02883_ keymem.key_mem\[6\]\[33\] _06010_ sky130_fd_sc_hd__mux2_2
XFILLER_0_203_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22095_ VGND VPWR _01760_ _06530_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_160_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_121_1157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_238_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21046_ VGND VPWR _01268_ _05973_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_195_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_226_472 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_92_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24805_ VGND VPWR VPWR VGND clk _01298_ reset_n keymem.key_mem\[6\]\[30\] sky130_fd_sc_hd__dfrtp_2
X_25785_ keymem.prev_key1_reg\[101\] clk _02278_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_134_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22997_ VGND VPWR VGND VPWR _06888_ keymem.prev_key1_reg\[50\] _06965_ _02227_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_243_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24736_ VGND VPWR VPWR VGND clk _01229_ reset_n keymem.key_mem\[7\]\[89\] sky130_fd_sc_hd__dfrtp_2
X_12750_ VGND VPWR VGND VPWR _08295_ _07665_ keymem.key_mem\[4\]\[58\] _08292_ _08294_
+ sky130_fd_sc_hd__a211o_2
X_21948_ VGND VPWR VPWR VGND _06449_ _04933_ keymem.key_mem\[3\]\[39\] _06453_ sky130_fd_sc_hd__mux2_2
XFILLER_0_55_1074 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_214_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11701_ VGND VPWR result[17] _07414_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_96_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12681_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[52\] _07918_ keymem.key_mem\[10\]\[52\]
+ _08193_ _08232_ sky130_fd_sc_hd__a22o_2
X_24667_ VGND VPWR VPWR VGND clk _01160_ reset_n keymem.key_mem\[7\]\[20\] sky130_fd_sc_hd__dfrtp_2
X_21879_ VGND VPWR _01659_ _06415_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14420_ VPWR VGND VPWR VGND _09889_ _09607_ _09888_ sky130_fd_sc_hd__or2_2
XFILLER_0_132_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11632_ VPWR VGND VGND VPWR _07372_ encdec next sky130_fd_sc_hd__nand2_2
X_23618_ VGND VPWR VPWR VGND clk _00119_ reset_n keymem.key_mem\[14\]\[107\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_166_265 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24598_ VGND VPWR VPWR VGND clk _01091_ reset_n keymem.key_mem\[8\]\[79\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_25_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14351_ VGND VPWR VPWR VGND _09178_ _09658_ _09821_ _09820_ _09819_ sky130_fd_sc_hd__o211a_2
XPHY_EDGE_ROW_95_2_Left_566 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23549_ VGND VPWR VPWR VGND clk _00050_ reset_n keymem.key_mem\[14\]\[38\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_53_948 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13302_ VPWR VGND VPWR VGND _08791_ keymem.key_mem\[5\]\[113\] _08052_ keymem.key_mem\[13\]\[113\]
+ _07695_ _08792_ sky130_fd_sc_hd__a221o_2
XFILLER_0_18_691 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17070_ VPWR VGND VPWR VGND _03190_ key[64] _08935_ sky130_fd_sc_hd__or2_2
X_14282_ VPWR VGND VGND VPWR _09751_ _09752_ _09747_ sky130_fd_sc_hd__nor2_2
X_16021_ _11339_ _11476_ _11338_ _11291_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_25219_ VGND VPWR VPWR VGND clk _01712_ reset_n keymem.key_mem\[3\]\[60\] sky130_fd_sc_hd__dfrtp_2
X_13233_ VPWR VGND VPWR VGND _08729_ keymem.key_mem\[11\]\[106\] _08011_ keymem.key_mem\[2\]\[106\]
+ _07733_ _08730_ sky130_fd_sc_hd__a221o_2
XFILLER_0_27_1154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13164_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[99\] _08577_ _08667_ _08663_ _08668_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_221_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12115_ VGND VPWR _07712_ _07711_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17972_ VGND VPWR _03577_ _03912_ _03913_ _03738_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_13095_ VGND VPWR enc_block.round_key\[92\] _08605_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19711_ VGND VPWR VPWR VGND _05259_ keymem.key_mem\[11\]\[16\] _11447_ _05263_ sky130_fd_sc_hd__mux2_2
XFILLER_0_100_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16923_ VGND VPWR VPWR VGND _02986_ keymem.key_mem\[14\]\[50\] _03056_ _03057_ sky130_fd_sc_hd__mux2_2
X_12046_ VGND VPWR _07646_ _07545_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_137_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_264_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_205_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19642_ VGND VPWR _00613_ _05224_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16854_ VGND VPWR VGND VPWR _09866_ key[172] _02994_ _02993_ sky130_fd_sc_hd__a21oi_2
X_15805_ VPWR VGND VPWR VGND _11192_ _11208_ _11197_ _11225_ _11261_ sky130_fd_sc_hd__or4_2
X_19573_ VPWR VGND keymem.key_mem\[12\]\[80\] _05189_ _05173_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13997_ VGND VPWR VGND VPWR _09320_ _09354_ _09468_ _09329_ _09373_ _09469_ sky130_fd_sc_hd__o32a_2
X_16785_ VGND VPWR VPWR VGND _09521_ key[166] keymem.prev_key1_reg\[38\] _02931_ sky130_fd_sc_hd__mux2_2
XFILLER_0_254_1388 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_38_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18524_ VGND VPWR _04403_ _04400_ _04402_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15736_ VGND VPWR VGND VPWR _11192_ _11191_ _11190_ keymem.prev_key1_reg\[22\] _08955_
+ _08942_ sky130_fd_sc_hd__a32o_2
X_12948_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[78\] _07771_ keymem.key_mem\[2\]\[78\]
+ _07546_ _08473_ sky130_fd_sc_hd__a22o_2
XFILLER_0_204_188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18455_ VGND VPWR _04340_ enc_block.block_w1_reg\[26\] enc_block.block_w1_reg\[31\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15667_ VGND VPWR VGND VPWR _10565_ _10513_ _10667_ _10511_ _11124_ sky130_fd_sc_hd__o22a_2
X_12879_ VPWR VGND VPWR VGND _08410_ keymem.key_mem\[11\]\[71\] _08090_ keymem.key_mem\[2\]\[71\]
+ _08131_ _08411_ sky130_fd_sc_hd__a221o_2
XFILLER_0_134_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17406_ VGND VPWR VGND VPWR _03489_ _02911_ keylen _03490_ sky130_fd_sc_hd__a21o_2
XFILLER_0_150_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14618_ VGND VPWR _10086_ _09868_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18386_ VPWR VGND VGND VPWR _04279_ _04024_ _04277_ sky130_fd_sc_hd__nand2_2
X_15598_ VGND VPWR _11056_ keymem.prev_key0_reg\[14\] _11055_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_263 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14549_ VPWR VGND VGND VPWR _10016_ _09651_ _09059_ _09230_ _09061_ _10017_ sky130_fd_sc_hd__a311o_2
X_17337_ VPWR VGND keymem.prev_key0_reg\[92\] _03429_ _02771_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_15_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_125_140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17268_ VGND VPWR VPWR VGND _02539_ _02540_ keymem.prev_key0_reg\[85\] _03367_ sky130_fd_sc_hd__or3_2
XFILLER_0_109_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_650 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19007_ VPWR VGND VPWR VGND _04836_ _04788_ _04835_ enc_block.block_w2_reg\[26\]
+ _04613_ _00366_ sky130_fd_sc_hd__a221o_2
X_16219_ VGND VPWR VPWR VGND _11567_ _11521_ _02383_ _02384_ sky130_fd_sc_hd__or3_2
XFILLER_0_24_672 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_52_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17199_ VPWR VGND VPWR VGND _03305_ _03303_ _03301_ key[205] _03027_ _03306_ sky130_fd_sc_hd__a221o_2
XFILLER_0_109_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_491 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_115_2_Right_187 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_80_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_355 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_87_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_545 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19909_ VGND VPWR _00738_ _05366_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_122_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_243_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22920_ VGND VPWR VGND VPWR _06918_ _02495_ _03860_ _06884_ _02548_ sky130_fd_sc_hd__a211o_2
XFILLER_0_194_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22851_ VPWR VGND VGND VPWR keymem.round_ctr_rst _05241_ _06873_ _02173_ sky130_fd_sc_hd__nor3_2
XFILLER_0_97_119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_194_1291 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_39_1058 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_116_1204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_998 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21802_ VGND VPWR _01625_ _06372_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25570_ VGND VPWR VPWR VGND clk _02063_ reset_n keymem.key_mem\[0\]\[27\] sky130_fd_sc_hd__dfrtp_2
X_22782_ VGND VPWR VPWR VGND _06784_ keymem.key_mem\[0\]\[90\] _03418_ _06852_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24521_ VGND VPWR VPWR VGND clk _01014_ reset_n keymem.key_mem\[8\]\[2\] sky130_fd_sc_hd__dfrtp_2
X_21733_ VGND VPWR VGND VPWR _06259_ _03226_ _01592_ _06336_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_148_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24452_ VGND VPWR VPWR VGND clk _00945_ reset_n keymem.key_mem\[9\]\[61\] sky130_fd_sc_hd__dfrtp_2
X_21664_ VGND VPWR _01559_ _06300_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_148_287 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_455 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_46_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23403_ VGND VPWR _07274_ enc_block.block_w0_reg\[19\] enc_block.block_w0_reg\[23\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20615_ VGND VPWR _01069_ _05741_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24383_ VGND VPWR VPWR VGND clk _00876_ reset_n keymem.key_mem\[10\]\[120\] sky130_fd_sc_hd__dfrtp_2
X_21595_ VGND VPWR _01526_ _06264_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_89_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_233 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23334_ VGND VPWR _07212_ enc_block.block_w0_reg\[21\] _07211_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20546_ VGND VPWR _01036_ _05705_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_127_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23265_ VGND VPWR _07150_ enc_block.block_w2_reg\[5\] _07149_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20477_ VGND VPWR VPWR VGND _05660_ _03627_ keymem.key_mem\[9\]\[121\] _05668_ sky130_fd_sc_hd__mux2_2
XFILLER_0_28_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25004_ VGND VPWR VPWR VGND clk _01497_ reset_n keymem.key_mem\[5\]\[101\] sky130_fd_sc_hd__dfrtp_2
X_22216_ VGND VPWR _01816_ _06595_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_161_1_Right_762 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23196_ VGND VPWR _07087_ enc_block.block_w2_reg\[7\] _07086_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22147_ VGND VPWR VPWR VGND _06554_ _10098_ keymem.key_mem\[2\]\[4\] _06559_ sky130_fd_sc_hd__mux2_2
XFILLER_0_30_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_140_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_218_247 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22078_ VGND VPWR _01752_ _06521_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_246_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_22_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13920_ VGND VPWR _09392_ _09391_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21029_ VGND VPWR VPWR VGND _05956_ _05079_ keymem.key_mem\[7\]\[122\] _05963_ sky130_fd_sc_hd__mux2_2
XFILLER_0_199_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_57_1114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_236_1030 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13851_ VGND VPWR _09323_ _09322_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_230_902 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_138_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25837_ VGND VPWR VPWR VGND clk _02330_ reset_n enc_block.block_w3_reg\[25\] sky130_fd_sc_hd__dfrtp_2
X_12802_ VGND VPWR enc_block.round_key\[63\] _08341_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_241_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_35_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13782_ VGND VPWR _09254_ _09253_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_39_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16570_ VPWR VGND _02728_ _02727_ keymem.prev_key0_reg\[122\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_25768_ keymem.prev_key1_reg\[84\] clk _02261_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_96_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15521_ VPWR VGND VGND VPWR _10543_ _10572_ _10980_ _10563_ _10867_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_57_517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12733_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[57\] _07691_ keymem.key_mem\[7\]\[57\]
+ _08016_ _08279_ sky130_fd_sc_hd__a22o_2
XFILLER_0_139_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_96_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24719_ VGND VPWR VPWR VGND clk _01212_ reset_n keymem.key_mem\[7\]\[72\] sky130_fd_sc_hd__dfrtp_2
X_25699_ keymem.prev_key1_reg\[15\] clk _02192_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_123_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18240_ VPWR VGND VGND VPWR _04146_ _04147_ enc_block.round_key\[111\] sky130_fd_sc_hd__nor2_2
X_15452_ VGND VPWR VGND VPWR _10838_ key[139] _10901_ _10902_ _10913_ _10912_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_249_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12664_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[50\] _08216_ keymem.key_mem\[7\]\[50\]
+ _07703_ _08217_ sky130_fd_sc_hd__a22o_2
XFILLER_0_139_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14403_ VPWR VGND VPWR VGND _09437_ _09478_ _09397_ _09472_ _09872_ sky130_fd_sc_hd__or4_2
X_15383_ VPWR VGND VPWR VGND _10726_ _10843_ _10841_ _10577_ _10844_ sky130_fd_sc_hd__or4_2
XFILLER_0_26_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18171_ VPWR VGND _04084_ _04083_ enc_block.round_key\[105\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_249_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_414 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12595_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[43\] _08145_ _08154_ _08149_ _08155_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_92_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_84 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14334_ VPWR VGND VGND VPWR _09071_ _09105_ _09646_ _09804_ sky130_fd_sc_hd__nor3_2
X_17122_ VGND VPWR _00081_ _03236_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_40_406 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_68_1276 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17053_ VGND VPWR _00074_ _03174_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_208_1143 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14265_ VPWR VGND VGND VPWR _09735_ _09733_ _09734_ sky130_fd_sc_hd__nand2_2
X_16004_ VPWR VGND VPWR VGND _11173_ _11248_ _11247_ _11233_ _11459_ sky130_fd_sc_hd__or4_2
XFILLER_0_46_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13216_ VGND VPWR _08714_ _07534_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14196_ VPWR VGND VGND VPWR _09667_ _09184_ _09666_ sky130_fd_sc_hd__nand2_2
XFILLER_0_20_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13147_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[98\] _07685_ keymem.key_mem\[2\]\[98\]
+ _07697_ _08652_ sky130_fd_sc_hd__a22o_2
XFILLER_0_209_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_57_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17955_ VGND VPWR _00249_ _03901_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13078_ VGND VPWR VGND VPWR _07841_ keymem.key_mem\[4\]\[91\] _08587_ _08589_ _08590_
+ _08480_ sky130_fd_sc_hd__a2111o_2
X_16906_ VGND VPWR VPWR VGND _03041_ keymem.prev_key1_reg\[81\] _11450_ _11451_ _08927_
+ sky130_fd_sc_hd__o31a_2
X_12029_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[2\] _07596_ keymem.key_mem\[12\]\[2\]
+ _07578_ _07630_ sky130_fd_sc_hd__a22o_2
XFILLER_0_228_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17886_ VGND VPWR _00227_ _03854_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_164_14 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_442 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19625_ VGND VPWR _00605_ _05215_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16837_ VPWR VGND VGND VPWR _02978_ _10903_ _10904_ sky130_fd_sc_hd__nand2_2
XFILLER_0_75_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_251_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19556_ VGND VPWR _00572_ _05179_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16768_ VGND VPWR VPWR VGND _09521_ key[165] keymem.prev_key1_reg\[37\] _02915_ sky130_fd_sc_hd__mux2_2
XFILLER_0_92_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_215_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18507_ VPWR VGND VPWR VGND _04387_ block[71] _03979_ enc_block.block_w0_reg\[7\]
+ _04138_ _04388_ sky130_fd_sc_hd__a221o_2
XFILLER_0_177_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15719_ enc_block.sword_ctr_reg\[1\] _11175_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[17\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_75_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19487_ VGND VPWR VPWR VGND _05138_ _04935_ keymem.key_mem\[12\]\[40\] _05143_ sky130_fd_sc_hd__mux2_2
XFILLER_0_48_539 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16699_ VGND VPWR VGND VPWR _02844_ _02843_ keymem.prev_key1_reg\[127\] _02852_ sky130_fd_sc_hd__a21o_2
X_18438_ _04323_ _04325_ _04294_ _04324_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_267_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_282 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_150_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_111_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_44_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_12_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18369_ VPWR VGND VPWR VGND _04263_ block[123] _03958_ enc_block.block_w0_reg\[27\]
+ _03953_ _04264_ sky130_fd_sc_hd__a221o_2
XFILLER_0_17_948 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20400_ VGND VPWR VPWR VGND _05627_ _03364_ keymem.key_mem\[9\]\[84\] _05628_ sky130_fd_sc_hd__mux2_2
XFILLER_0_160_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21380_ VGND VPWR VPWR VGND _06140_ _02838_ keymem.key_mem\[5\]\[30\] _06150_ sky130_fd_sc_hd__mux2_2
XFILLER_0_82_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20331_ VGND VPWR VPWR VGND _05591_ _03068_ keymem.key_mem\[9\]\[51\] _05592_ sky130_fd_sc_hd__mux2_2
XFILLER_0_3_363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_305 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_98_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23050_ VGND VPWR VPWR VGND _02248_ _06996_ _03250_ _06976_ _06997_ sky130_fd_sc_hd__o31a_2
X_20262_ VGND VPWR _00902_ _05555_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_12_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22001_ VPWR VGND keymem.key_mem\[3\]\[64\] _06481_ _06469_ VPWR VGND sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_116_2_Right_188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20193_ VGND VPWR _00871_ _05517_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_23_Left_291 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_256_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_122_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1041 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_228_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_23_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_138_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23952_ VGND VPWR VPWR VGND clk _00445_ reset_n keymem.key_mem\[13\]\[73\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_196_1397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22903_ VGND VPWR VGND VPWR _02191_ _06907_ _06882_ keymem.prev_key1_reg\[14\] sky130_fd_sc_hd__o21a_2
XFILLER_0_157_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_212_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23883_ VGND VPWR VPWR VGND clk _00376_ reset_n keymem.key_mem\[13\]\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25622_ VGND VPWR VPWR VGND clk _02115_ reset_n keymem.key_mem\[0\]\[79\] sky130_fd_sc_hd__dfrtp_2
X_22834_ VPWR VGND VGND VPWR _06865_ keymem.rcon_reg\[0\] keymem.rcon_logic.tmp_rcon\[0\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_195_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25553_ VGND VPWR VPWR VGND clk _02046_ reset_n keymem.key_mem\[0\]\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22765_ VGND VPWR _02115_ _06845_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24504_ VGND VPWR VPWR VGND clk _00997_ reset_n keymem.key_mem\[9\]\[113\] sky130_fd_sc_hd__dfrtp_2
X_21716_ VGND VPWR _01584_ _06327_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_176_360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25484_ VGND VPWR VPWR VGND clk _01977_ reset_n keymem.key_mem\[1\]\[69\] sky130_fd_sc_hd__dfrtp_2
X_22696_ VGND VPWR _02073_ _06818_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_93_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_712 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24435_ VGND VPWR VPWR VGND clk _00928_ reset_n keymem.key_mem\[9\]\[44\] sky130_fd_sc_hd__dfrtp_2
X_21647_ VGND VPWR _01551_ _06291_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_30_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24366_ VGND VPWR VPWR VGND clk _00859_ reset_n keymem.key_mem\[10\]\[103\] sky130_fd_sc_hd__dfrtp_2
X_12380_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[24\] _07649_ keymem.key_mem\[2\]\[24\]
+ _07697_ _07959_ sky130_fd_sc_hd__a22o_2
XFILLER_0_164_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21578_ VGND VPWR _01520_ _06253_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_168_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_78_2_Right_150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23317_ VPWR VGND VGND VPWR _07196_ _07197_ _07194_ sky130_fd_sc_hd__nor2_2
XFILLER_0_104_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20529_ VGND VPWR _01028_ _05696_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24297_ VGND VPWR VPWR VGND clk _00790_ reset_n keymem.key_mem\[10\]\[34\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_166_1190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_158_1_Left_425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14050_ VGND VPWR _09522_ _09521_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23248_ _07133_ _07135_ _03955_ _07134_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_13001_ VGND VPWR VGND VPWR _08521_ _08150_ keymem.key_mem\[3\]\[83\] _08518_ _08520_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_249_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_162_1_Right_763 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23179_ VPWR VGND VGND VPWR _07076_ _03929_ _06892_ sky130_fd_sc_hd__nand2_2
XFILLER_0_101_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_140_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_101_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17740_ VGND VPWR _00177_ _03758_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14952_ VGND VPWR VGND VPWR _10416_ enc_block.sword_ctr_reg\[0\] enc_block.block_w1_reg\[12\]
+ enc_block.sword_ctr_reg\[1\] sky130_fd_sc_hd__and3b_2
XFILLER_0_265_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13903_ VGND VPWR _09375_ _09374_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_175_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17671_ VGND VPWR _00156_ _03710_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14883_ VPWR VGND VPWR VGND _09042_ _10347_ _09181_ _09840_ _10348_ sky130_fd_sc_hd__a22o_2
XFILLER_0_242_570 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19410_ VPWR VGND keymem.key_mem\[12\]\[5\] _05101_ _05095_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16622_ VPWR VGND VPWR VGND _02778_ keymem.prev_key1_reg\[92\] sky130_fd_sc_hd__inv_2
X_13834_ VGND VPWR _09306_ _09275_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_43_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19341_ VGND VPWR VPWR VGND _05046_ _05054_ keymem.key_mem\[13\]\[110\] _05055_ sky130_fd_sc_hd__mux2_2
X_13765_ VPWR VGND VPWR VGND _09227_ _09236_ _09233_ _09220_ _09237_ sky130_fd_sc_hd__or4_2
X_16553_ VGND VPWR VGND VPWR _02710_ _02709_ _02711_ _02712_ sky130_fd_sc_hd__a21o_2
XFILLER_0_169_1208 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15504_ VPWR VGND VGND VPWR _10735_ _10916_ _10963_ _10964_ sky130_fd_sc_hd__nor3_2
XFILLER_0_84_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12716_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[55\] _07748_ keymem.key_mem\[4\]\[55\]
+ _07734_ _08264_ sky130_fd_sc_hd__a22o_2
X_19272_ VPWR VGND keymem.key_mem_we _05010_ _03383_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13696_ VGND VPWR _09168_ _09077_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_112_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16484_ VGND VPWR VGND VPWR _02644_ _02643_ _02645_ keymem.prev_key0_reg\[23\] sky130_fd_sc_hd__a21oi_2
XFILLER_0_26_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18223_ VPWR VGND VGND VPWR _04130_ _04131_ _03966_ sky130_fd_sc_hd__nor2_2
X_15435_ VPWR VGND _10896_ keymem.prev_key0_reg\[75\] keymem.prev_key0_reg\[43\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
X_12647_ VGND VPWR enc_block.round_key\[48\] _08201_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_112_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_26_745 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_186_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_182_374 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18154_ VPWR VGND VGND VPWR _04068_ _03983_ _04067_ sky130_fd_sc_hd__nand2_2
X_15366_ VPWR VGND _10828_ _10827_ keymem.prev_key1_reg\[106\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_12578_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[42\] _07649_ keymem.key_mem\[11\]\[42\]
+ _07658_ _08139_ sky130_fd_sc_hd__a22o_2
XFILLER_0_182_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17105_ VPWR VGND _10077_ _03221_ _10078_ VPWR VGND sky130_fd_sc_hd__and2_2
X_14317_ VGND VPWR VGND VPWR _09786_ _09785_ _09787_ _09784_ _09566_ sky130_fd_sc_hd__nand4_2
XFILLER_0_83_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15297_ VGND VPWR VGND VPWR _10759_ _10758_ _10703_ _10670_ _10548_ sky130_fd_sc_hd__and4_2
X_18085_ VPWR VGND VGND VPWR _04005_ _04004_ _10827_ sky130_fd_sc_hd__nand2_2
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17036_ VPWR VGND VPWR VGND _03159_ key[189] _10322_ sky130_fd_sc_hd__or2_2
X_14248_ VGND VPWR _09719_ _08935_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_22_973 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_223_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_150_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_878 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14179_ VGND VPWR VGND VPWR _09649_ _09648_ _09650_ _09647_ _09645_ sky130_fd_sc_hd__nand4_2
XFILLER_0_237_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18987_ VPWR VGND VPWR VGND _04818_ block[56] _04744_ enc_block.block_w2_reg\[24\]
+ _04798_ _04819_ sky130_fd_sc_hd__a221o_2
XFILLER_0_84_11 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_193_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17938_ VGND VPWR VPWR VGND _03874_ _03889_ keymem.prev_key0_reg\[103\] _03890_ sky130_fd_sc_hd__mux2_2
XFILLER_0_175_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_193_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17869_ VGND VPWR VPWR VGND _03836_ _03842_ keymem.prev_key0_reg\[81\] _03843_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_172_2_Left_643 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_261_890 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19608_ VGND VPWR VPWR VGND _05205_ _05027_ keymem.key_mem\[12\]\[97\] _05207_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20880_ VGND VPWR VGND VPWR _05884_ keymem.key_mem_we _03068_ _05864_ _01191_ sky130_fd_sc_hd__a31o_2
XFILLER_0_205_294 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_49_804 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19539_ VGND VPWR VGND VPWR _05170_ keymem.key_mem_we _03194_ _05164_ _00564_ sky130_fd_sc_hd__a31o_2
XFILLER_0_220_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_152_1278 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22550_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[76\] _06754_ _06753_ _04992_ _01984_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_75_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_130_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21501_ VGND VPWR _01483_ _06213_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_723 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22481_ VGND VPWR VPWR VGND _06726_ keymem.key_mem\[1\]\[35\] _02904_ _06734_ sky130_fd_sc_hd__mux2_2
XFILLER_0_9_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_734 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_12_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24220_ VGND VPWR VPWR VGND clk _00713_ reset_n keymem.key_mem\[11\]\[85\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_133_216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21432_ VGND VPWR _01450_ _06177_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_90_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24151_ VGND VPWR VPWR VGND clk _00644_ reset_n keymem.key_mem\[11\]\[16\] sky130_fd_sc_hd__dfrtp_2
X_21363_ VGND VPWR _01417_ _06141_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_86_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23102_ VGND VPWR VGND VPWR _03438_ _03437_ _03442_ _07028_ sky130_fd_sc_hd__a21o_2
X_20314_ VGND VPWR VPWR VGND _05580_ _02985_ keymem.key_mem\[9\]\[43\] _05583_ sky130_fd_sc_hd__mux2_2
X_24082_ VGND VPWR VPWR VGND clk _00575_ reset_n keymem.key_mem\[12\]\[75\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_101_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21294_ VGND VPWR _01386_ _06103_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_241_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23033_ VGND VPWR VGND VPWR _06986_ _03204_ _03860_ _03208_ _06951_ sky130_fd_sc_hd__a211o_2
X_20245_ VGND VPWR VPWR VGND _05546_ _10836_ keymem.key_mem\[9\]\[10\] _05547_ sky130_fd_sc_hd__mux2_2
XFILLER_0_198_1415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_2_Right_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_239_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20176_ VGND VPWR _00863_ _05508_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24984_ VGND VPWR VPWR VGND clk _01477_ reset_n keymem.key_mem\[5\]\[81\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_157_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23935_ VGND VPWR VPWR VGND clk _00428_ reset_n keymem.key_mem\[13\]\[56\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_235_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_224_592 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_197_934 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11880_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[11\] dec_new_block\[107\]
+ _07504_ sky130_fd_sc_hd__mux2_2
X_23866_ VGND VPWR VPWR VGND clk _00359_ reset_n enc_block.block_w2_reg\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25605_ VGND VPWR VPWR VGND clk _02098_ reset_n keymem.key_mem\[0\]\[62\] sky130_fd_sc_hd__dfrtp_2
X_22817_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[116\] _06860_ _06859_ _05066_ _02152_
+ sky130_fd_sc_hd__a22o_2
X_23797_ VGND VPWR VPWR VGND clk _00290_ reset_n enc_block.block_w0_reg\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_251_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_319 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13550_ VGND VPWR _09022_ _09021_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_55_807 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25536_ VGND VPWR VPWR VGND clk _02029_ reset_n keymem.key_mem\[1\]\[121\] sky130_fd_sc_hd__dfrtp_2
X_22748_ VPWR VGND VGND VPWR _06840_ keymem.key_mem\[0\]\[68\] _06839_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_11_Right_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_55_818 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_149_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12501_ VGND VPWR _08069_ _07746_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13481_ VPWR VGND VPWR VGND _08953_ enc_block.block_w0_reg\[2\] _08952_ sky130_fd_sc_hd__or2_2
X_25467_ VGND VPWR VPWR VGND clk _01960_ reset_n keymem.key_mem\[1\]\[52\] sky130_fd_sc_hd__dfrtp_2
X_22679_ VGND VPWR _02063_ _06811_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15220_ VGND VPWR VGND VPWR _10682_ _10639_ _10541_ _10644_ _10683_ sky130_fd_sc_hd__o22a_2
XFILLER_0_81_136 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24418_ VGND VPWR VPWR VGND clk _00911_ reset_n keymem.key_mem\[9\]\[27\] sky130_fd_sc_hd__dfrtp_2
X_12432_ VPWR VGND VPWR VGND _08005_ keymem.key_mem\[9\]\[29\] _07717_ keymem.key_mem\[10\]\[29\]
+ _07909_ _08006_ sky130_fd_sc_hd__a221o_2
X_25398_ VGND VPWR VPWR VGND clk _01891_ reset_n keymem.key_mem\[2\]\[111\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_129_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15151_ VGND VPWR VGND VPWR _10476_ _10538_ _10566_ _10569_ _10615_ sky130_fd_sc_hd__o22a_2
XFILLER_0_2_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12363_ VGND VPWR enc_block.round_key\[22\] _07943_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24349_ VGND VPWR VPWR VGND clk _00842_ reset_n keymem.key_mem\[10\]\[86\] sky130_fd_sc_hd__dfrtp_2
X_14102_ VGND VPWR VGND VPWR _09573_ _09309_ _09339_ _09328_ _09338_ sky130_fd_sc_hd__and4_2
XPHY_EDGE_ROW_79_2_Right_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_205_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15082_ VGND VPWR _10546_ _10545_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_65_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12294_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[17\] _07618_ keymem.key_mem\[12\]\[17\]
+ _07673_ _07880_ sky130_fd_sc_hd__a22o_2
XFILLER_0_146_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_267_949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14033_ VGND VPWR VGND VPWR _09455_ _09504_ _09505_ _09438_ _09471_ sky130_fd_sc_hd__nor4_2
X_18910_ VPWR VGND VPWR VGND _04749_ block[48] _04744_ enc_block.block_w3_reg\[16\]
+ _04666_ _04750_ sky130_fd_sc_hd__a221o_2
XFILLER_0_200_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_20_Right_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19890_ VGND VPWR _00729_ _05356_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18841_ VPWR VGND VPWR VGND _04687_ block[41] _03979_ enc_block.block_w0_reg\[9\]
+ _04138_ _04688_ sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_163_1_Right_764 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_105_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_684 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18772_ VGND VPWR _04625_ enc_block.block_w2_reg\[26\] _04624_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_1017 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15984_ VGND VPWR VPWR VGND keymem.round_ctr_reg\[0\] _11439_ _10653_ _11440_ sky130_fd_sc_hd__mux2_2
X_17723_ VGND VPWR VGND VPWR _03748_ keymem.prev_key0_reg\[29\] _00170_ _03736_ sky130_fd_sc_hd__a21bo_2
X_14935_ VGND VPWR VGND VPWR _10399_ enc_block.block_w2_reg\[10\] enc_block.sword_ctr_reg\[1\]
+ enc_block.sword_ctr_reg\[0\] sky130_fd_sc_hd__and3b_2
XFILLER_0_76_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_101_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_222_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_89_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_175_1278 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_89_247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_76_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17654_ VGND VPWR VPWR VGND _03681_ _03698_ keymem.prev_key0_reg\[10\] _03699_ sky130_fd_sc_hd__mux2_2
XFILLER_0_37_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14866_ VGND VPWR VGND VPWR _09141_ _09109_ _10331_ _09221_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_89_269 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_72_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16605_ VPWR VGND VPWR VGND _02762_ key[155] _10286_ sky130_fd_sc_hd__or2_2
X_13817_ VPWR VGND VPWR VGND _09289_ enc_block.block_w0_reg\[28\] _08995_ sky130_fd_sc_hd__or2_2
X_17585_ VPWR VGND VPWR VGND _03645_ key[252] _09927_ sky130_fd_sc_hd__or2_2
X_14797_ VGND VPWR VPWR VGND _10230_ _10262_ keymem.prev_key0_reg\[102\] _10263_ sky130_fd_sc_hd__or3_2
XFILLER_0_161_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19324_ VPWR VGND keymem.key_mem_we _05043_ _03525_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16536_ VGND VPWR VGND VPWR _09629_ _09589_ _02695_ _10360_ sky130_fd_sc_hd__a21oi_2
X_13748_ VPWR VGND VGND VPWR _09219_ _09218_ _09106_ _09059_ _09215_ _09220_ sky130_fd_sc_hd__a311o_2
XFILLER_0_112_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19255_ VPWR VGND keymem.key_mem\[13\]\[79\] _05000_ _04979_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16467_ VGND VPWR VGND VPWR _11235_ _11330_ _11336_ _11385_ _02628_ sky130_fd_sc_hd__o22a_2
X_13679_ VGND VPWR VGND VPWR _09138_ _09132_ _09116_ _09102_ _09151_ sky130_fd_sc_hd__o22a_2
X_18206_ VPWR VGND VPWR VGND _04116_ _03970_ _10961_ sky130_fd_sc_hd__or2_2
XFILLER_0_112_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15418_ VPWR VGND VPWR VGND _10879_ _10603_ _10635_ sky130_fd_sc_hd__or2_2
X_19186_ VPWR VGND keymem.key_mem_we _04958_ _03075_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16398_ VGND VPWR VGND VPWR _02559_ _11367_ _02560_ _11211_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_60_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1374 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_87_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_147_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18137_ VPWR VGND VGND VPWR _04052_ _04053_ _04041_ sky130_fd_sc_hd__nor2_2
X_15349_ VGND VPWR VPWR VGND _10478_ _10476_ _10580_ _10811_ sky130_fd_sc_hd__or3_2
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_748 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_83_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_388 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_48_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18068_ _03987_ _03989_ _03982_ _03988_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_83_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17019_ VGND VPWR _09931_ key[60] _03143_ _10327_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_229_139 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20030_ VGND VPWR VPWR VGND _05424_ _02934_ keymem.key_mem\[10\]\[38\] _05432_ sky130_fd_sc_hd__mux2_2
XFILLER_0_95_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_123_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21981_ VGND VPWR VGND VPWR _06470_ keymem.key_mem_we _03091_ _06446_ _01706_ sky130_fd_sc_hd__a31o_2
XFILLER_0_154_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_158_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23720_ keymem.prev_key0_reg\[76\] clk _00217_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_94_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20932_ VGND VPWR _05912_ _05819_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_55_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_359 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_7_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23651_ keymem.prev_key0_reg\[7\] clk _00148_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20863_ VGND VPWR _01183_ _05875_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_49_634 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_117_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_280 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22602_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[112\] _06777_ _06776_ _05058_ _02020_
+ sky130_fd_sc_hd__a22o_2
X_23582_ VGND VPWR VPWR VGND clk _00083_ reset_n keymem.key_mem\[14\]\[71\] sky130_fd_sc_hd__dfrtp_2
X_20794_ VGND VPWR _05838_ _05820_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25321_ VGND VPWR VPWR VGND clk _01814_ reset_n keymem.key_mem\[2\]\[34\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_130_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22533_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[66\] _06754_ _06753_ _04977_ _01974_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_63_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_146_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_108 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_130_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25252_ VGND VPWR VPWR VGND clk _01745_ reset_n keymem.key_mem\[3\]\[93\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_165_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22464_ VGND VPWR _06726_ _06701_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_267_1173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24203_ VGND VPWR VPWR VGND clk _00696_ reset_n keymem.key_mem\[11\]\[68\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_263_1037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21415_ VGND VPWR _01442_ _06168_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_165_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25183_ VGND VPWR VPWR VGND clk _01676_ reset_n keymem.key_mem\[3\]\[24\] sky130_fd_sc_hd__dfrtp_2
X_22395_ VGND VPWR VPWR VGND _06680_ _03633_ keymem.key_mem\[2\]\[122\] _06689_ sky130_fd_sc_hd__mux2_2
XFILLER_0_66_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_121_219 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_556 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24134_ VGND VPWR VPWR VGND clk _00627_ reset_n keymem.key_mem\[12\]\[127\] sky130_fd_sc_hd__dfrtp_2
X_21346_ VGND VPWR _01409_ _06132_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_245_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_898 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_205_Right_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24065_ VGND VPWR VPWR VGND clk _00558_ reset_n keymem.key_mem\[12\]\[58\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_206_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_163_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21277_ VGND VPWR _01378_ _06094_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_229_640 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23016_ VPWR VGND VGND VPWR _06977_ _03124_ _06976_ sky130_fd_sc_hd__nand2_2
X_20228_ VGND VPWR VPWR VGND _05535_ _09862_ keymem.key_mem\[9\]\[2\] _05538_ sky130_fd_sc_hd__mux2_2
XFILLER_0_229_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_102_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_246_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_835 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_141_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1220 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_244_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20159_ VGND VPWR _00855_ _05499_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_102_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_805 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_176_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12981_ VGND VPWR VGND VPWR _08503_ _07665_ keymem.key_mem\[4\]\[81\] _08500_ _08502_
+ sky130_fd_sc_hd__a211o_2
X_24967_ VGND VPWR VPWR VGND clk _01460_ reset_n keymem.key_mem\[5\]\[64\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_172_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_1001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_73_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14720_ VPWR VGND _10187_ _10186_ keymem.prev_key0_reg\[101\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_231_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23918_ VGND VPWR VPWR VGND clk _00411_ reset_n keymem.key_mem\[13\]\[39\] sky130_fd_sc_hd__dfrtp_2
X_11932_ VGND VPWR _07535_ _07534_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24898_ VGND VPWR VPWR VGND clk _01391_ reset_n keymem.key_mem\[6\]\[123\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_214_Right_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_73_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_764 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11863_ VGND VPWR result[98] _07495_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14651_ VGND VPWR VPWR VGND _09398_ _09348_ _09247_ _10118_ sky130_fd_sc_hd__or3_2
X_23849_ VGND VPWR VPWR VGND clk _00342_ reset_n enc_block.block_w2_reg\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_213_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13602_ VPWR VGND VPWR VGND _09063_ _09073_ _09070_ _09056_ _09074_ sky130_fd_sc_hd__or4_2
X_17370_ VPWR VGND VPWR VGND _03458_ _02677_ _03456_ key[223] _10838_ _03459_ sky130_fd_sc_hd__a221o_2
X_14582_ VPWR VGND VGND VPWR _09419_ _10050_ _09349_ sky130_fd_sc_hd__nor2_2
X_11794_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[0\] dec_new_block\[64\]
+ _07461_ sky130_fd_sc_hd__mux2_2
XFILLER_0_27_306 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16321_ VPWR VGND VPWR VGND _02484_ keymem.prev_key1_reg\[85\] sky130_fd_sc_hd__inv_2
X_13533_ VGND VPWR _09005_ _09004_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_113_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25519_ VGND VPWR VPWR VGND clk _02012_ reset_n keymem.key_mem\[1\]\[104\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_211_1172 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_10_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19040_ VGND VPWR _04866_ enc_block.round_key\[62\] _04865_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_16252_ VPWR VGND VGND VPWR _02416_ _02414_ _02415_ sky130_fd_sc_hd__nand2_2
XFILLER_0_183_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13464_ VGND VPWR _08936_ _08935_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_42_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15203_ VPWR VGND _09679_ _10666_ _09708_ VPWR VGND sky130_fd_sc_hd__and2_2
X_12415_ VPWR VGND VPWR VGND _07990_ keymem.key_mem\[11\]\[27\] _07600_ keymem.key_mem\[10\]\[27\]
+ _07561_ _07991_ sky130_fd_sc_hd__a221o_2
XFILLER_0_183_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16183_ VGND VPWR VPWR VGND _11477_ _11262_ _11376_ _02348_ sky130_fd_sc_hd__or3_2
X_13395_ VGND VPWR enc_block.round_key\[122\] _08875_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_223_Right_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15134_ VPWR VGND VGND VPWR _10496_ _10598_ _10565_ sky130_fd_sc_hd__nor2_2
XFILLER_0_224_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12346_ VGND VPWR VGND VPWR _07924_ keymem.key_mem\[9\]\[21\] _07925_ _07927_ _07928_
+ _07616_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_23_578 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15065_ VGND VPWR VPWR VGND _10403_ _10466_ _10439_ _10529_ sky130_fd_sc_hd__or3_2
XFILLER_0_267_746 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_224_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19942_ VGND VPWR _00754_ _05383_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12277_ VGND VPWR VGND VPWR _07753_ keymem.key_mem\[8\]\[16\] _07860_ _07863_ _07864_
+ _07616_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_10_239 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_49_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14016_ VGND VPWR VGND VPWR _09330_ _09268_ _09312_ _09487_ _09488_ sky130_fd_sc_hd__o22a_2
X_19873_ VGND VPWR _00721_ _05347_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_177_1307 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_120_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18824_ VPWR VGND _04673_ _04672_ enc_block.round_key\[39\] VPWR VGND sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_164_1_Right_765 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_120_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_65_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18755_ _04608_ _04610_ _04560_ _04609_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_15967_ VGND VPWR VGND VPWR _11329_ _11313_ _11327_ _11422_ _11222_ _11423_ sky130_fd_sc_hd__o32a_2
XFILLER_0_190_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_890 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17706_ VGND VPWR _03736_ _03729_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_164_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_236_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14918_ VGND VPWR VGND VPWR _10381_ _10371_ _10372_ _10377_ _10382_ sky130_fd_sc_hd__a31o_2
X_18686_ VPWR VGND VPWR VGND _04547_ block[90] _04487_ enc_block.block_w1_reg\[26\]
+ _04543_ _04548_ sky130_fd_sc_hd__a221o_2
X_15898_ VPWR VGND VPWR VGND _11350_ _11353_ _11354_ _11346_ _11347_ sky130_fd_sc_hd__or4b_2
XFILLER_0_76_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17637_ VGND VPWR VPWR VGND _03679_ key[133] keymem.prev_key1_reg\[5\] _03687_ sky130_fd_sc_hd__mux2_2
X_14849_ VPWR VGND VGND VPWR _09457_ _09585_ _10313_ _10314_ sky130_fd_sc_hd__nor3_2
XFILLER_0_37_1167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_33_1009 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_231_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_370 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_105_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_965 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_187_285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17568_ VGND VPWR VGND VPWR _02728_ _02342_ _03630_ _03629_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_105_63 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_45_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19307_ VGND VPWR VPWR VGND _05025_ _05031_ keymem.key_mem\[13\]\[99\] _05032_ sky130_fd_sc_hd__mux2_2
X_16519_ VGND VPWR keymem.prev_key1_reg\[120\] _02668_ _02679_ _02669_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_18_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17499_ VGND VPWR _02866_ key[113] _03570_ _10189_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_19238_ VGND VPWR VGND VPWR _04988_ keymem.key_mem_we _03268_ _04968_ _00445_ sky130_fd_sc_hd__a31o_2
XFILLER_0_6_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19169_ VPWR VGND keymem.key_mem_we _04947_ _03015_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_26_394 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_48_1230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21200_ VGND VPWR _01341_ _06054_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_197_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_170_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22180_ VGND VPWR _01799_ _06576_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_147_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_48_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21131_ VGND VPWR _06018_ _05971_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_2_973 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_69_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_223_1054 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21062_ VGND VPWR _01276_ _05981_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_195_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20013_ VGND VPWR VPWR VGND _05413_ _02839_ keymem.key_mem\[10\]\[30\] _05423_ sky130_fd_sc_hd__mux2_2
X_24821_ VGND VPWR VPWR VGND clk _01314_ reset_n keymem.key_mem\[6\]\[46\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_236_1415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_198_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_119_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_55_1212 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21964_ VPWR VGND keymem.key_mem\[3\]\[47\] _06461_ _06439_ VPWR VGND sky130_fd_sc_hd__and2_2
X_24752_ VGND VPWR VPWR VGND clk _01245_ reset_n keymem.key_mem\[7\]\[105\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_94_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20915_ VGND VPWR VGND VPWR _05903_ keymem.key_mem_we _03217_ _05893_ _01207_ sky130_fd_sc_hd__a31o_2
X_23703_ keymem.prev_key0_reg\[59\] clk _00200_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_222_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24683_ VGND VPWR VPWR VGND clk _01176_ reset_n keymem.key_mem\[7\]\[36\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_6_Left_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21895_ VPWR VGND keymem.key_mem\[3\]\[15\] _06424_ _06413_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_16_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_167_1_Left_434 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_55_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23634_ VGND VPWR VPWR VGND clk _00135_ reset_n keymem.key_mem\[14\]\[123\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_138_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20846_ VGND VPWR VGND VPWR _05866_ keymem.key_mem_we _02904_ _05864_ _01175_ sky130_fd_sc_hd__a31o_2
XFILLER_0_230_1047 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_2_Left_606 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_64_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23565_ VGND VPWR VPWR VGND clk _00066_ reset_n keymem.key_mem\[14\]\[54\] sky130_fd_sc_hd__dfrtp_2
X_20777_ VPWR VGND keymem.key_mem\[7\]\[4\] _05829_ _05824_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_9_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_851 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22516_ VGND VPWR _01966_ _06745_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25304_ VGND VPWR VPWR VGND clk _01797_ reset_n keymem.key_mem\[2\]\[17\] sky130_fd_sc_hd__dfrtp_2
X_23496_ VPWR VGND VPWR VGND _07356_ _03950_ _07355_ enc_block.block_w3_reg\[30\]
+ _07126_ _02335_ sky130_fd_sc_hd__a221o_2
XFILLER_0_52_629 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1038 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_134_355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25235_ VGND VPWR VPWR VGND clk _01728_ reset_n keymem.key_mem\[3\]\[76\] sky130_fd_sc_hd__dfrtp_2
X_22447_ VGND VPWR _01925_ _06717_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_165_1244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_165_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12200_ VGND VPWR _07793_ _07644_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_66_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13180_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[101\] _08216_ keymem.key_mem\[2\]\[101\]
+ _08131_ _08682_ sky130_fd_sc_hd__a22o_2
X_25166_ VGND VPWR VPWR VGND clk _01659_ reset_n keymem.key_mem\[3\]\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22378_ VGND VPWR _06680_ _06552_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_241_1121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_249_724 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12131_ VGND VPWR VGND VPWR _07728_ _07721_ keymem.key_mem\[14\]\[6\] _07723_ _07727_
+ sky130_fd_sc_hd__a211o_2
X_24117_ VGND VPWR VPWR VGND clk _00610_ reset_n keymem.key_mem\[12\]\[110\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_248_223 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21329_ VGND VPWR _01401_ _06123_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_27_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25097_ VGND VPWR VPWR VGND clk _01590_ reset_n keymem.key_mem\[4\]\[66\] sky130_fd_sc_hd__dfrtp_2
X_24048_ VGND VPWR VPWR VGND clk _00541_ reset_n keymem.key_mem\[12\]\[41\] sky130_fd_sc_hd__dfrtp_2
X_12062_ VGND VPWR _07662_ _07572_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_102_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16870_ VPWR VGND VGND VPWR _02947_ _11055_ _11092_ _03008_ sky130_fd_sc_hd__nor3_2
XFILLER_0_198_1086 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_205_805 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15821_ VPWR VGND VPWR VGND _11268_ _11276_ _11271_ _11260_ _11277_ sky130_fd_sc_hd__or4_2
XFILLER_0_245_996 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_176_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_99_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18540_ VGND VPWR _04417_ _04354_ _04416_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_137_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15752_ VGND VPWR VGND VPWR _11208_ _11201_ _11200_ keymem.prev_key1_reg\[21\] _10402_
+ _09255_ sky130_fd_sc_hd__a32o_2
XFILLER_0_38_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_176_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12964_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[80\] _07568_ keymem.key_mem\[6\]\[80\]
+ _07759_ _08487_ sky130_fd_sc_hd__a22o_2
XFILLER_0_73_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_1_Left_366 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14703_ _09185_ _10170_ _09047_ _09945_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_137_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11915_ VGND VPWR result[124] _07521_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18471_ VPWR VGND _04355_ enc_block.block_w1_reg\[28\] enc_block.block_w2_reg\[20\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_15683_ VPWR VGND VGND VPWR _10789_ _11139_ _10939_ _10719_ _11140_ sky130_fd_sc_hd__and4b_2
XPHY_EDGE_ROW_67_2_Left_538 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_73_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1272 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12895_ VPWR VGND VPWR VGND _08424_ keymem.key_mem\[1\]\[73\] _07715_ keymem.key_mem\[2\]\[73\]
+ _07546_ _08425_ sky130_fd_sc_hd__a221o_2
XFILLER_0_200_510 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_34_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17422_ VGND VPWR VPWR VGND _09730_ _03503_ key[230] _03504_ sky130_fd_sc_hd__mux2_2
X_14634_ VPWR VGND _10101_ keymem.prev_key1_reg\[37\] keymem.prev_key1_reg\[5\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
X_11846_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[26\] dec_new_block\[90\]
+ _07487_ sky130_fd_sc_hd__mux2_2
XFILLER_0_51_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17353_ VGND VPWR _03444_ _03443_ VPWR VGND sky130_fd_sc_hd__buf_1
X_11777_ VGND VPWR result[55] _07452_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14565_ VPWR VGND VGND VPWR _09437_ _09466_ _10033_ _09302_ _09444_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_136 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_55_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_222_50 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16304_ VGND VPWR VPWR VGND _02468_ _10386_ _02465_ _02466_ _02467_ sky130_fd_sc_hd__o31a_2
X_13516_ VPWR VGND VPWR VGND _08988_ enc_block.block_w0_reg\[5\] _08952_ sky130_fd_sc_hd__or2_2
XFILLER_0_55_478 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17284_ VGND VPWR VGND VPWR _03381_ _03380_ _03382_ keylen sky130_fd_sc_hd__a21oi_2
X_14496_ VGND VPWR VGND VPWR _09961_ _09189_ _09962_ _09963_ _09965_ _09964_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_183_1311 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_148_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19023_ VPWR VGND VPWR VGND _04850_ block[60] _04837_ enc_block.block_w2_reg\[28\]
+ _04798_ _04851_ sky130_fd_sc_hd__a221o_2
XFILLER_0_187_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16235_ VPWR VGND _02400_ _02399_ keymem.prev_key0_reg\[19\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_152_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_125_366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13447_ VGND VPWR _08922_ _08921_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_10_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_320 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_109_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_148_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16166_ _10775_ _11620_ _07386_ _10814_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_13378_ VPWR VGND VPWR VGND _08859_ keymem.key_mem\[14\]\[121\] _08032_ keymem.key_mem\[4\]\[121\]
+ _07637_ _08860_ sky130_fd_sc_hd__a221o_2
XFILLER_0_144_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_181_2_Left_652 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_258 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15117_ VGND VPWR VGND VPWR _10581_ _10580_ _10579_ _10578_ sky130_fd_sc_hd__o21a_2
X_12329_ VGND VPWR _07912_ _07600_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_45_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16097_ VGND VPWR VGND VPWR _11551_ _11550_ _11549_ _09521_ sky130_fd_sc_hd__o21a_2
X_15048_ VPWR VGND VGND VPWR _10511_ _10512_ _10508_ sky130_fd_sc_hd__nor2_2
X_19925_ VGND VPWR VPWR VGND _05372_ keymem.key_mem\[11\]\[118\] _03607_ _05375_ sky130_fd_sc_hd__mux2_2
XFILLER_0_255_738 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_259_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19856_ VGND VPWR _00713_ _05338_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_236_963 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_263_760 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_165_1_Right_766 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18807_ VGND VPWR _04657_ enc_block.block_w2_reg\[29\] enc_block.block_w0_reg\[14\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_19787_ VGND VPWR _00680_ _05302_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_194_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16999_ _02735_ _03125_ _03124_ _02736_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_250_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_155_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18738_ VPWR VGND VGND VPWR _04594_ _04591_ _04593_ sky130_fd_sc_hd__nand2_2
XFILLER_0_56_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_91_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_155_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18669_ VPWR VGND VPWR VGND _04532_ block[88] _04487_ enc_block.block_w1_reg\[24\]
+ _04425_ _04533_ sky130_fd_sc_hd__a221o_2
XFILLER_0_116_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1323 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_8_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20700_ VGND VPWR VPWR VGND _05783_ _03480_ keymem.key_mem\[8\]\[98\] _05786_ sky130_fd_sc_hd__mux2_2
XFILLER_0_153_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21680_ VGND VPWR VPWR VGND _06308_ _02985_ keymem.key_mem\[4\]\[43\] _06309_ sky130_fd_sc_hd__mux2_2
XFILLER_0_8_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20631_ VGND VPWR VPWR VGND _05747_ _03202_ keymem.key_mem\[8\]\[65\] _05750_ sky130_fd_sc_hd__mux2_2
XFILLER_0_231_1389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_175_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1255 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_116_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23350_ VPWR VGND VPWR VGND _07226_ block[14] _03980_ enc_block.block_w1_reg\[14\]
+ _03978_ _07227_ sky130_fd_sc_hd__a221o_2
XFILLER_0_50_1186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20562_ VGND VPWR _01044_ _05713_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_15_821 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22301_ VGND VPWR VPWR VGND _06634_ _03306_ keymem.key_mem\[2\]\[77\] _06640_ sky130_fd_sc_hd__mux2_2
XFILLER_0_166_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23281_ VPWR VGND VGND VPWR _07126_ _07165_ _04062_ sky130_fd_sc_hd__nor2_2
XFILLER_0_127_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20493_ VGND VPWR VPWR VGND _05676_ _09536_ keymem.key_mem\[8\]\[0\] _05677_ sky130_fd_sc_hd__mux2_2
XFILLER_0_26_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25020_ VGND VPWR VPWR VGND clk _01513_ reset_n keymem.key_mem\[5\]\[117\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_166_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22232_ VGND VPWR VPWR VGND _06600_ _02998_ keymem.key_mem\[2\]\[44\] _06604_ sky130_fd_sc_hd__mux2_2
XFILLER_0_30_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1082 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_242_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22163_ VPWR VGND VGND VPWR _06568_ keymem.key_mem\[2\]\[11\] _06567_ sky130_fd_sc_hd__nand2_2
XFILLER_0_24_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21114_ VGND VPWR _01300_ _06009_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22094_ VGND VPWR VPWR VGND _06527_ _05050_ keymem.key_mem\[3\]\[108\] _06530_ sky130_fd_sc_hd__mux2_2
XFILLER_0_258_598 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_203_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21045_ VGND VPWR VPWR VGND _05972_ _09536_ keymem.key_mem\[6\]\[0\] _05973_ sky130_fd_sc_hd__mux2_2
XFILLER_0_201_1160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_91 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_253_270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_236_1223 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24804_ VGND VPWR VPWR VGND clk _01297_ reset_n keymem.key_mem\[6\]\[29\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_173_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25784_ keymem.prev_key1_reg\[100\] clk _02277_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22996_ VGND VPWR VPWR VGND _03050_ _03048_ _06965_ _06881_ _03054_ sky130_fd_sc_hd__o211a_2
XFILLER_0_232_1109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24735_ VGND VPWR VPWR VGND clk _01228_ reset_n keymem.key_mem\[7\]\[88\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_214_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_178 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21947_ VGND VPWR _01690_ _06452_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_96_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11700_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[17\] dec_new_block\[17\]
+ _07414_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12680_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[52\] _07652_ keymem.key_mem\[6\]\[52\]
+ _07657_ _08231_ sky130_fd_sc_hd__a22o_2
XFILLER_0_214_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_913 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21878_ VGND VPWR VPWR VGND _06403_ _04889_ keymem.key_mem\[3\]\[7\] _06415_ sky130_fd_sc_hd__mux2_2
X_24666_ VGND VPWR VPWR VGND clk _01159_ reset_n keymem.key_mem\[7\]\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_96_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_210_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11631_ VGND VPWR VGND VPWR _00005_ aes_core_ctrl_reg\[0\] next aes_core_ctrl_reg\[1\]
+ _07371_ _07366_ sky130_fd_sc_hd__a32o_2
X_20829_ VGND VPWR VGND VPWR _05857_ keymem.key_mem_we _02765_ _05850_ _01167_ sky130_fd_sc_hd__a31o_2
X_23617_ VGND VPWR VPWR VGND clk _00118_ reset_n keymem.key_mem\[14\]\[106\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24597_ VGND VPWR VPWR VGND clk _01090_ reset_n keymem.key_mem\[8\]\[78\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_166_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_181_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14350_ VGND VPWR VGND VPWR _09019_ _09149_ _09103_ _09196_ _09058_ _09820_ sky130_fd_sc_hd__o32a_2
XFILLER_0_64_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_64_264 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23548_ VGND VPWR VPWR VGND clk _00049_ reset_n keymem.key_mem\[14\]\[37\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_107_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_110_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13301_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[113\] _07651_ keymem.key_mem\[6\]\[113\]
+ _07656_ _08791_ sky130_fd_sc_hd__a22o_2
X_14281_ VGND VPWR VGND VPWR _09751_ _09748_ _09419_ _09341_ _09750_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_24_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_437 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23479_ VGND VPWR VGND VPWR _07341_ _04149_ _07093_ _07342_ enc_block.block_w3_reg\[28\]
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_134_163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16020_ VPWR VGND VPWR VGND _11472_ _11474_ _11475_ _11463_ _11468_ sky130_fd_sc_hd__or4b_2
X_13232_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[106\] _07742_ keymem.key_mem\[8\]\[106\]
+ _07903_ _08729_ sky130_fd_sc_hd__a22o_2
X_25218_ VGND VPWR VPWR VGND clk _01711_ reset_n keymem.key_mem\[3\]\[59\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_492 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13163_ VGND VPWR VGND VPWR _08667_ _07877_ keymem.key_mem\[10\]\[99\] _08664_ _08666_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_0_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25149_ VGND VPWR VPWR VGND clk _01642_ reset_n keymem.key_mem\[4\]\[118\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_1166 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_221_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12114_ VGND VPWR _07711_ _07565_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_206_1093 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17971_ VPWR VGND VPWR VGND _03912_ keymem.prev_key1_reg\[114\] sky130_fd_sc_hd__inv_2
X_13094_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[92\] _08577_ _08604_ _08600_ _08605_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_221_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19710_ VGND VPWR _00643_ _05262_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16922_ VGND VPWR VGND VPWR _03056_ _03054_ _03050_ _03048_ _03055_ sky130_fd_sc_hd__o211ai_2
X_12045_ VGND VPWR _07645_ _07644_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_46_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_900 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19641_ VGND VPWR VPWR VGND _05216_ _05060_ keymem.key_mem\[12\]\[113\] _05224_ sky130_fd_sc_hd__mux2_2
XFILLER_0_205_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16853_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[76\] keymem.prev_key1_reg\[44\]
+ _02993_ _02992_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_233_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_232_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15804_ VPWR VGND VGND VPWR _11259_ _11260_ _11257_ sky130_fd_sc_hd__nor2_2
X_19572_ VGND VPWR VGND VPWR _05188_ keymem.key_mem_we _03322_ _05187_ _00579_ sky130_fd_sc_hd__a31o_2
X_16784_ VPWR VGND VPWR VGND _02930_ keymem.prev_key1_reg\[38\] sky130_fd_sc_hd__inv_2
X_13996_ VPWR VGND VGND VPWR _09247_ _09468_ _09447_ sky130_fd_sc_hd__nor2_2
X_18523_ VPWR VGND _04402_ _04401_ _04319_ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_153_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15735_ VPWR VGND VPWR VGND _11191_ enc_block.block_w0_reg\[22\] _09273_ sky130_fd_sc_hd__or2_2
XFILLER_0_204_178 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12947_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[78\] _07588_ keymem.key_mem\[14\]\[78\]
+ _07984_ _08472_ sky130_fd_sc_hd__a22o_2
XFILLER_0_38_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18454_ VPWR VGND VPWR VGND _04339_ _04291_ _04338_ enc_block.block_w1_reg\[2\] _04317_
+ _00310_ sky130_fd_sc_hd__a221o_2
X_15666_ VGND VPWR VGND VPWR _10608_ _10575_ _10543_ _10639_ _11123_ sky130_fd_sc_hd__o22a_2
XFILLER_0_5_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12878_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[71\] _07667_ keymem.key_mem\[8\]\[71\]
+ _07540_ _08410_ sky130_fd_sc_hd__a22o_2
XFILLER_0_56_710 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_8_807 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17405_ VPWR VGND VGND VPWR _03489_ key[228] _10967_ sky130_fd_sc_hd__nand2_2
X_14617_ VGND VPWR _10085_ _09722_ VPWR VGND sky130_fd_sc_hd__buf_1
X_11829_ VGND VPWR result[81] _07478_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18385_ VPWR VGND VPWR VGND _04278_ _04024_ _04277_ sky130_fd_sc_hd__or2_2
XFILLER_0_5_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15597_ VPWR VGND _11055_ keymem.prev_key0_reg\[78\] keymem.prev_key0_reg\[46\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_150_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_328 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17336_ VGND VPWR _00103_ _03428_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_185_1417 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14548_ VGND VPWR VGND VPWR _09052_ _09072_ _10016_ _09007_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_102_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17267_ VGND VPWR _03366_ _09543_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_125_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14479_ VGND VPWR VGND VPWR _09948_ _09050_ _09140_ _09099_ _09167_ _09105_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_70_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_226_1425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_523 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19006_ VPWR VGND VGND VPWR _04778_ _04836_ _04256_ sky130_fd_sc_hd__nor2_2
XFILLER_0_109_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16218_ VGND VPWR VGND VPWR _11390_ _11266_ _11280_ _11210_ _02383_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_30_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_23_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17198_ VGND VPWR VGND VPWR _03304_ _11034_ _03305_ keylen sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_49_Right_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_52_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_109_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_578 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16149_ VGND VPWR VGND VPWR _11236_ _11336_ _11205_ _11320_ _11603_ sky130_fd_sc_hd__o22a_2
XFILLER_0_23_194 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_178_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_367 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_87_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_11_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1046 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_209_930 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19908_ VGND VPWR VPWR VGND _05361_ keymem.key_mem\[11\]\[110\] _03555_ _05366_ sky130_fd_sc_hd__mux2_2
XFILLER_0_194_56 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19839_ VGND VPWR VPWR VGND _05328_ keymem.key_mem\[11\]\[77\] _03306_ _05330_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_166_1_Right_767 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_224_966 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22850_ VGND VPWR VGND VPWR keymem.round_ctr_reg\[0\] keymem.key_mem_we _06873_ keymem.round_ctr_reg\[1\]
+ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_58_Right_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_78_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_251_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_190_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_116_1216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21801_ VGND VPWR VPWR VGND _06366_ _03499_ keymem.key_mem\[4\]\[101\] _06372_ sky130_fd_sc_hd__mux2_2
XFILLER_0_116_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22781_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[89\] _06850_ _06849_ _05015_ _02125_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_17_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21732_ VPWR VGND VGND VPWR _06259_ _06336_ keymem.key_mem\[4\]\[68\] sky130_fd_sc_hd__nor2_2
X_24520_ VGND VPWR VPWR VGND clk _01013_ reset_n keymem.key_mem\[8\]\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1248 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_233 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24451_ VGND VPWR VPWR VGND clk _00944_ reset_n keymem.key_mem\[9\]\[60\] sky130_fd_sc_hd__dfrtp_2
X_21663_ VGND VPWR VPWR VGND _06297_ _02903_ keymem.key_mem\[4\]\[35\] _06300_ sky130_fd_sc_hd__mux2_2
XFILLER_0_231_1186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_143_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23402_ VPWR VGND VPWR VGND _07273_ _04874_ _07272_ enc_block.block_w3_reg\[19\]
+ _07126_ _02324_ sky130_fd_sc_hd__a221o_2
X_20614_ VGND VPWR VPWR VGND _05736_ _03118_ keymem.key_mem\[8\]\[57\] _05741_ sky130_fd_sc_hd__mux2_2
XFILLER_0_163_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_46_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24382_ VGND VPWR VPWR VGND clk _00875_ reset_n keymem.key_mem\[10\]\[119\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_163_236 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21594_ VGND VPWR VPWR VGND _06263_ _09861_ keymem.key_mem\[4\]\[2\] _06264_ sky130_fd_sc_hd__mux2_2
XFILLER_0_7_862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23333_ VPWR VGND _07211_ enc_block.block_w1_reg\[12\] enc_block.block_w3_reg\[29\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_116_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_89_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20545_ VGND VPWR VPWR VGND _05703_ _02688_ keymem.key_mem\[8\]\[24\] _05705_ sky130_fd_sc_hd__mux2_2
XFILLER_0_62_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_50_919 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_127_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23264_ VGND VPWR _07149_ enc_block.block_w3_reg\[29\] enc_block.block_w1_reg\[14\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20476_ VGND VPWR _01004_ _05667_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_67_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25003_ VGND VPWR VPWR VGND clk _01496_ reset_n keymem.key_mem\[5\]\[100\] sky130_fd_sc_hd__dfrtp_2
X_22215_ VGND VPWR VPWR VGND _06589_ _02913_ keymem.key_mem\[2\]\[36\] _06595_ sky130_fd_sc_hd__mux2_2
XFILLER_0_28_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23195_ VPWR VGND _07086_ enc_block.block_w3_reg\[31\] enc_block.block_w3_reg\[24\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_24_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22146_ VGND VPWR _01783_ _06558_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_98_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22077_ VGND VPWR VPWR VGND _06516_ _05033_ keymem.key_mem\[3\]\[100\] _06521_ sky130_fd_sc_hd__mux2_2
X_21028_ VGND VPWR _01261_ _05962_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_22_1085 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_261_538 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_227_793 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_254_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13850_ VPWR VGND VPWR VGND _09307_ _09309_ _09321_ _09275_ _09322_ sky130_fd_sc_hd__or4_2
X_25836_ VGND VPWR VPWR VGND clk _02329_ reset_n enc_block.block_w3_reg\[24\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1332 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12801_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[63\] _07645_ _08340_ _08336_ _08341_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_199_678 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_74_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13781_ VGND VPWR VGND VPWR _09253_ _09252_ _09002_ keymem.prev_key1_reg\[27\] _09003_
+ _09251_ sky130_fd_sc_hd__a32o_2
X_25767_ keymem.prev_key1_reg\[83\] clk _02260_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_35_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22979_ VGND VPWR VGND VPWR _06955_ _02977_ _06891_ _02984_ _06951_ sky130_fd_sc_hd__a211o_2
XFILLER_0_198_188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15520_ VPWR VGND VPWR VGND _10979_ keymem.prev_key0_reg\[109\] sky130_fd_sc_hd__inv_2
X_24718_ VGND VPWR VPWR VGND clk _01211_ reset_n keymem.key_mem\[7\]\[71\] sky130_fd_sc_hd__dfrtp_2
X_12732_ VGND VPWR enc_block.round_key\[56\] _08278_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_35_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25698_ keymem.prev_key1_reg\[14\] clk _02191_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_214_1384 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15451_ VPWR VGND VPWR VGND _10909_ _10908_ _10912_ _10911_ keylen sky130_fd_sc_hd__a211oi_2
XFILLER_0_96_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_38_743 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12663_ VGND VPWR _08216_ _07618_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24649_ VGND VPWR VPWR VGND clk _01142_ reset_n keymem.key_mem\[7\]\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_249_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_916 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14402_ VGND VPWR VPWR VGND _09871_ _09338_ _09307_ _09285_ _09336_ sky130_fd_sc_hd__o31a_2
X_18170_ VPWR VGND VPWR VGND _04082_ block[105] _04076_ enc_block.block_w2_reg\[9\]
+ _04007_ _04083_ sky130_fd_sc_hd__a221o_2
X_15382_ VGND VPWR _10842_ _10547_ _10843_ _10644_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_12594_ VGND VPWR VGND VPWR _08154_ _08150_ keymem.key_mem\[3\]\[43\] _08151_ _08153_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_25_426 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_949 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_249_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17121_ VGND VPWR VPWR VGND _03185_ keymem.key_mem\[14\]\[69\] _03235_ _03236_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_25_437 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14333_ VPWR VGND VGND VPWR _09132_ _09803_ _09108_ sky130_fd_sc_hd__nor2_2
XFILLER_0_92_392 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17052_ VGND VPWR VPWR VGND _03084_ keymem.key_mem\[14\]\[62\] _03173_ _03174_ sky130_fd_sc_hd__mux2_2
XFILLER_0_145_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14264_ VGND VPWR VGND VPWR _09323_ _09388_ _09440_ _09565_ _09734_ sky130_fd_sc_hd__o22a_2
XFILLER_0_122_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_243_1046 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16003_ VGND VPWR VGND VPWR _10728_ _10677_ _11458_ keymem.round_ctr_reg\[0\] sky130_fd_sc_hd__a21oi_2
XFILLER_0_106_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13215_ VGND VPWR enc_block.round_key\[104\] _08713_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_204_1019 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_46_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14195_ VGND VPWR VGND VPWR _09666_ _09005_ _09045_ _09014_ _09001_ sky130_fd_sc_hd__and4_2
XFILLER_0_122_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1079 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13146_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[98\] _07834_ keymem.key_mem\[7\]\[98\]
+ _07650_ _08651_ sky130_fd_sc_hd__a22o_2
XFILLER_0_148_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_264_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17954_ VGND VPWR VPWR VGND _03896_ _03900_ keymem.prev_key0_reg\[108\] _03901_ sky130_fd_sc_hd__mux2_2
X_13077_ VPWR VGND VPWR VGND _08588_ keymem.key_mem\[10\]\[91\] _07909_ keymem.key_mem\[1\]\[91\]
+ _07715_ _08589_ sky130_fd_sc_hd__a221o_2
XFILLER_0_265_866 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_264_354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_178_1254 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16905_ VGND VPWR keymem.prev_key1_reg\[81\] _11450_ _03040_ _11451_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_256_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12028_ VGND VPWR _07629_ _07561_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17885_ VGND VPWR VPWR VGND _03836_ _03853_ keymem.prev_key0_reg\[86\] _03854_ sky130_fd_sc_hd__mux2_2
XFILLER_0_205_410 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_206_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16836_ VGND VPWR VPWR VGND _02977_ _10735_ _02974_ _02975_ _02976_ sky130_fd_sc_hd__o31a_2
X_19624_ VGND VPWR VPWR VGND _05205_ _05043_ keymem.key_mem\[12\]\[105\] _05215_ sky130_fd_sc_hd__mux2_2
XFILLER_0_79_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_117_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_156_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19555_ VGND VPWR VPWR VGND _05151_ _04986_ keymem.key_mem\[12\]\[72\] _05179_ sky130_fd_sc_hd__mux2_2
X_16767_ VGND VPWR _00048_ _02914_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13979_ VGND VPWR VPWR VGND _09444_ _09451_ _09353_ _09383_ _09450_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_53_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1070 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18506_ VPWR VGND VGND VPWR _04386_ _04387_ _04382_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_90_1_Right_691 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15718_ VGND VPWR _11174_ _11173_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_244_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19486_ VGND VPWR _00539_ _05142_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16698_ VGND VPWR VPWR VGND _11109_ _02850_ key[31] _02851_ sky130_fd_sc_hd__mux2_2
X_18437_ VPWR VGND VGND VPWR _04324_ _04318_ _04322_ sky130_fd_sc_hd__nand2_2
X_15649_ VPWR VGND VGND VPWR _11106_ keymem.prev_key1_reg\[79\] _11105_ sky130_fd_sc_hd__nand2_2
XFILLER_0_267_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18368_ _04261_ _04263_ _04064_ _04262_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_51_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_111_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_724 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_267_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17319_ VPWR VGND VGND VPWR _03412_ _03413_ keylen sky130_fd_sc_hd__nor2_2
XFILLER_0_32_908 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18299_ VGND VPWR VGND VPWR _02458_ _02430_ _04073_ _04201_ sky130_fd_sc_hd__a21o_2
XFILLER_0_44_779 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20330_ VGND VPWR _05591_ _05534_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_31_429 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_82_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_124_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20261_ VGND VPWR VPWR VGND _05546_ _02340_ keymem.key_mem\[9\]\[18\] _05555_ sky130_fd_sc_hd__mux2_2
XFILLER_0_3_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22000_ VGND VPWR VGND VPWR _06480_ keymem.key_mem_we _03184_ _06475_ _01715_ sky130_fd_sc_hd__a31o_2
XFILLER_0_12_676 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_256_822 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_204_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20192_ VGND VPWR VPWR VGND _05515_ _03585_ keymem.key_mem\[10\]\[115\] _05517_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_176_1_Left_443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_855 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_122_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_144_2_Left_615 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_243_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23951_ VGND VPWR VPWR VGND clk _00444_ reset_n keymem.key_mem\[13\]\[72\] sky130_fd_sc_hd__dfrtp_2
X_22902_ VGND VPWR VGND VPWR _06907_ _11054_ _03860_ _06884_ _11097_ sky130_fd_sc_hd__a211o_2
X_23882_ VGND VPWR VPWR VGND clk _00375_ reset_n keymem.key_mem\[13\]\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_212_914 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_212_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_167_1_Right_768 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_93_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25621_ VGND VPWR VPWR VGND clk _02114_ reset_n keymem.key_mem\[0\]\[78\] sky130_fd_sc_hd__dfrtp_2
X_22833_ VPWR VGND keymem.key_mem_we _06864_ _06861_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_17_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25552_ VGND VPWR VPWR VGND clk _02045_ reset_n keymem.key_mem\[0\]\[9\] sky130_fd_sc_hd__dfrtp_2
X_22764_ VGND VPWR VPWR VGND _06833_ keymem.key_mem\[0\]\[79\] _03322_ _06845_ sky130_fd_sc_hd__mux2_2
XFILLER_0_211_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24503_ VGND VPWR VPWR VGND clk _00996_ reset_n keymem.key_mem\[9\]\[112\] sky130_fd_sc_hd__dfrtp_2
X_21715_ VGND VPWR VPWR VGND _06319_ _03149_ keymem.key_mem\[4\]\[60\] _06327_ sky130_fd_sc_hd__mux2_2
X_22695_ VGND VPWR VPWR VGND _06809_ keymem.key_mem\[0\]\[37\] _02924_ _06818_ sky130_fd_sc_hd__mux2_2
X_25483_ VGND VPWR VPWR VGND clk _01976_ reset_n keymem.key_mem\[1\]\[68\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_47_551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_52_1089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_176_383 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24434_ VGND VPWR VPWR VGND clk _00927_ reset_n keymem.key_mem\[9\]\[43\] sky130_fd_sc_hd__dfrtp_2
X_21646_ VGND VPWR VPWR VGND _06286_ _02764_ keymem.key_mem\[4\]\[27\] _06291_ sky130_fd_sc_hd__mux2_2
XFILLER_0_93_178 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_30_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24365_ VGND VPWR VPWR VGND clk _00858_ reset_n keymem.key_mem\[10\]\[102\] sky130_fd_sc_hd__dfrtp_2
X_21577_ VGND VPWR VPWR VGND _06116_ _03647_ keymem.key_mem\[5\]\[124\] _06253_ sky130_fd_sc_hd__mux2_2
XFILLER_0_23_908 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23316_ VGND VPWR _07196_ _07118_ _07195_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20528_ VGND VPWR VPWR VGND _05692_ _11446_ keymem.key_mem\[8\]\[16\] _05696_ sky130_fd_sc_hd__mux2_2
X_24296_ VGND VPWR VPWR VGND clk _00789_ reset_n keymem.key_mem\[10\]\[33\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_104_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_249_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23247_ VPWR VGND VPWR VGND _07134_ _07128_ _07132_ sky130_fd_sc_hd__or2_2
X_20459_ VGND VPWR _00996_ _05658_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_28_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13000_ VPWR VGND VPWR VGND _08519_ keymem.key_mem\[14\]\[83\] _07706_ keymem.key_mem\[4\]\[83\]
+ _07854_ _08520_ sky130_fd_sc_hd__a221o_2
XFILLER_0_24_1125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_682 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23178_ VGND VPWR _02298_ _07075_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_76_2_Left_547 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_140_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_238_Left_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_247_866 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22129_ VGND VPWR VPWR VGND _06538_ _05085_ keymem.key_mem\[3\]\[125\] _06548_ sky130_fd_sc_hd__mux2_2
XFILLER_0_262_803 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_140_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14951_ enc_block.sword_ctr_reg\[1\] _10415_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[12\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_101_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13902_ VPWR VGND VPWR VGND _09328_ _09309_ _09285_ _09338_ _09374_ sky130_fd_sc_hd__or4_2
X_17670_ VGND VPWR VPWR VGND _03703_ _03709_ keymem.prev_key0_reg\[15\] _03710_ sky130_fd_sc_hd__mux2_2
XFILLER_0_199_431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14882_ VGND VPWR VGND VPWR _10346_ _09190_ _09114_ _09057_ _10347_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_215_763 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_261_379 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16621_ VGND VPWR VGND VPWR _02768_ _02767_ keymem.prev_key1_reg\[124\] _02777_ sky130_fd_sc_hd__a21o_2
X_13833_ VGND VPWR VGND VPWR _09305_ _09246_ _09300_ _09303_ _09304_ sky130_fd_sc_hd__a211o_2
X_25819_ VGND VPWR VPWR VGND clk _02312_ reset_n enc_block.block_w3_reg\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_134_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19340_ VPWR VGND keymem.key_mem_we _05054_ _03555_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16552_ VPWR VGND VPWR VGND _02711_ keymem.prev_key1_reg\[89\] sky130_fd_sc_hd__inv_2
X_13764_ VPWR VGND VGND VPWR _09235_ _09234_ _09047_ _09041_ _09061_ _09236_ sky130_fd_sc_hd__a311o_2
XFILLER_0_134_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_468 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_190_2_Left_661 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_70_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15503_ VGND VPWR _10963_ keymem.prev_key0_reg\[108\] _10962_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_247_Left_514 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12715_ VGND VPWR VGND VPWR _07786_ keymem.key_mem\[10\]\[55\] _08260_ _08262_ _08263_
+ _08243_ sky130_fd_sc_hd__a2111o_2
X_19271_ VGND VPWR _00457_ _05009_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16483_ VGND VPWR VGND VPWR _02642_ _02640_ _02644_ _02641_ sky130_fd_sc_hd__nand3_2
XFILLER_0_214_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_151_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13695_ VGND VPWR _09167_ _09166_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_167_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18222_ VGND VPWR _04130_ _04127_ _04129_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_127_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15434_ VGND VPWR keymem.prev_key0_reg\[107\] _10839_ _10895_ _10893_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_26_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_84_178 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12646_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[48\] _08145_ _08200_ _08196_ _08201_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_84_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_53_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_249_1266 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_210_1089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18153_ VGND VPWR _04067_ enc_block.block_w2_reg\[15\] _04066_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_129_1_Right_730 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15365_ VPWR VGND VGND VPWR _10827_ _09827_ _09850_ sky130_fd_sc_hd__nand2_2
XFILLER_0_53_554 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12577_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[42\] _07690_ keymem.key_mem\[6\]\[42\]
+ _08137_ _08138_ sky130_fd_sc_hd__a22o_2
X_17104_ VGND VPWR VPWR VGND _10371_ _10089_ _03219_ _03220_ sky130_fd_sc_hd__mux2_2
X_14316_ VGND VPWR VGND VPWR _09466_ _09456_ _09450_ _09786_ sky130_fd_sc_hd__a21o_2
X_18084_ VGND VPWR _04004_ _03972_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_1285 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15296_ VPWR VGND VGND VPWR _10629_ _10482_ _10644_ _10547_ _10758_ _10757_ sky130_fd_sc_hd__o221a_2
XFILLER_0_25_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_802 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17035_ _02803_ _03158_ _03156_ _02804_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_14247_ VGND VPWR VGND VPWR _09717_ _09715_ _09713_ _09714_ _09718_ sky130_fd_sc_hd__a31o_2
XFILLER_0_262_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_264_Right_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_180_1166 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_256_Left_523 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14178_ VGND VPWR VGND VPWR _09646_ _09099_ _09007_ _09053_ _09649_ sky130_fd_sc_hd__o22a_2
XFILLER_0_0_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13129_ VGND VPWR VGND VPWR _08050_ keymem.key_mem\[7\]\[96\] _08633_ _08635_ _08636_
+ _07896_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_239_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_194_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18986_ _04816_ _04818_ _04560_ _04817_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_225_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_23 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17937_ VGND VPWR VGND VPWR _03508_ keymem.prev_key1_reg\[103\] _03889_ _03818_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_193_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_108_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17868_ VGND VPWR _03337_ _11449_ _03842_ _03789_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_117_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19607_ VGND VPWR _00596_ _05206_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16819_ VGND VPWR VGND VPWR _10740_ _10739_ _02962_ _02961_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_220_210 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_191_1262 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17799_ VGND VPWR VGND VPWR _03124_ _03792_ _03795_ _03793_ _03727_ _03796_ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_18_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_265_Left_532 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_49_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19538_ VPWR VGND keymem.key_mem\[12\]\[64\] _05170_ _05158_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_191_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_1_Right_692 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_165_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_18_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19469_ VGND VPWR VPWR VGND _05092_ _04920_ keymem.key_mem\[12\]\[32\] _05133_ sky130_fd_sc_hd__mux2_2
XFILLER_0_9_935 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_359 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_192_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21500_ VGND VPWR VPWR VGND _06209_ _03392_ keymem.key_mem\[5\]\[87\] _06213_ sky130_fd_sc_hd__mux2_2
XFILLER_0_130_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22480_ VGND VPWR _01942_ _06733_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_173_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_63_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_1027 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21431_ VGND VPWR VPWR VGND _06173_ _03090_ keymem.key_mem\[5\]\[54\] _06177_ sky130_fd_sc_hd__mux2_2
XFILLER_0_99_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24150_ VGND VPWR VPWR VGND clk _00643_ reset_n keymem.key_mem\[11\]\[15\] sky130_fd_sc_hd__dfrtp_2
X_21362_ VGND VPWR VPWR VGND _06140_ _02549_ keymem.key_mem\[5\]\[21\] _06141_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_640 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_31_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20313_ VGND VPWR _00926_ _05582_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23101_ VGND VPWR _02269_ _07027_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_31_248 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24081_ VGND VPWR VPWR VGND clk _00574_ reset_n keymem.key_mem\[12\]\[74\] sky130_fd_sc_hd__dfrtp_2
X_21293_ VGND VPWR VPWR VGND _06098_ _03607_ keymem.key_mem\[6\]\[118\] _06103_ sky130_fd_sc_hd__mux2_2
XFILLER_0_25_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_226_1085 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23032_ VGND VPWR VGND VPWR _02242_ _06985_ _06954_ keymem.prev_key1_reg\[65\] sky130_fd_sc_hd__o21a_2
XPHY_EDGE_ROW_231_Right_100 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20244_ VGND VPWR _05546_ _05534_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_40_793 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_99_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20175_ VGND VPWR VPWR VGND _05504_ _03538_ keymem.key_mem\[10\]\[107\] _05508_ sky130_fd_sc_hd__mux2_2
XFILLER_0_239_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24983_ VGND VPWR VPWR VGND clk _01476_ reset_n keymem.key_mem\[5\]\[80\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_239_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23934_ VGND VPWR VPWR VGND clk _00427_ reset_n keymem.key_mem\[13\]\[55\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_157_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23865_ VGND VPWR VPWR VGND clk _00358_ reset_n enc_block.block_w2_reg\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_168_103 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_168_1_Right_769 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25604_ VGND VPWR VPWR VGND clk _02097_ reset_n keymem.key_mem\[0\]\[61\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_36_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22816_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[115\] _06860_ _06859_ _05064_ _02151_
+ sky130_fd_sc_hd__a22o_2
X_23796_ VGND VPWR VPWR VGND clk _00289_ reset_n enc_block.block_w0_reg\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_66_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_251_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25535_ VGND VPWR VPWR VGND clk _02028_ reset_n keymem.key_mem\[1\]\[120\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_489 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_183_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22747_ VGND VPWR _06839_ _06784_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_109_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12500_ VPWR VGND VPWR VGND _08067_ keymem.key_mem\[14\]\[35\] _08003_ keymem.key_mem\[8\]\[35\]
+ _07655_ _08068_ sky130_fd_sc_hd__a221o_2
XFILLER_0_183_139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13480_ VGND VPWR _08952_ _08951_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25466_ VGND VPWR VPWR VGND clk _01959_ reset_n keymem.key_mem\[1\]\[51\] sky130_fd_sc_hd__dfrtp_2
X_22678_ VGND VPWR VPWR VGND _06809_ keymem.key_mem\[0\]\[27\] _02765_ _06811_ sky130_fd_sc_hd__mux2_2
XFILLER_0_63_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24417_ VGND VPWR VPWR VGND clk _00910_ reset_n keymem.key_mem\[9\]\[26\] sky130_fd_sc_hd__dfrtp_2
X_12431_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[29\] _07659_ keymem.key_mem\[6\]\[29\]
+ _07639_ _08005_ sky130_fd_sc_hd__a22o_2
XFILLER_0_168_1253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21629_ VGND VPWR VPWR VGND _06275_ _02409_ keymem.key_mem\[4\]\[19\] _06282_ sky130_fd_sc_hd__mux2_2
XFILLER_0_30_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_340 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25397_ VGND VPWR VPWR VGND clk _01890_ reset_n keymem.key_mem\[2\]\[110\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15150_ VGND VPWR VGND VPWR _10455_ _10565_ _10612_ _10614_ sky130_fd_sc_hd__a21o_2
XFILLER_0_50_513 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24348_ VGND VPWR VPWR VGND clk _00841_ reset_n keymem.key_mem\[10\]\[85\] sky130_fd_sc_hd__dfrtp_2
X_12362_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[22\] _07535_ _07942_ _07938_ _07943_
+ sky130_fd_sc_hd__o22a_2
X_14101_ VPWR VGND VGND VPWR _09366_ _09572_ _09318_ sky130_fd_sc_hd__nor2_2
X_15081_ VGND VPWR _10545_ _10544_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12293_ VPWR VGND VPWR VGND keymem.key_mem\[8\]\[17\] _07878_ keymem.key_mem\[4\]\[17\]
+ _07734_ _07879_ sky130_fd_sc_hd__a22o_2
XFILLER_0_50_568 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_107_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24279_ VGND VPWR VPWR VGND clk _00772_ reset_n keymem.key_mem\[10\]\[16\] sky130_fd_sc_hd__dfrtp_2
X_14032_ VPWR VGND VPWR VGND _09492_ _09503_ _09497_ _09483_ _09504_ sky130_fd_sc_hd__or4_2
XFILLER_0_82_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_247_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18840_ VPWR VGND VGND VPWR _04686_ _04687_ _03965_ sky130_fd_sc_hd__nor2_2
XFILLER_0_257_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18771_ VGND VPWR _04624_ enc_block.block_w2_reg\[31\] enc_block.block_w0_reg\[11\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15983_ VPWR VGND _11301_ _11439_ _11438_ VPWR VGND sky130_fd_sc_hd__and2_2
X_17722_ VGND VPWR VPWR VGND _03729_ _03747_ _02808_ _03748_ sky130_fd_sc_hd__or3_2
X_14934_ enc_block.sword_ctr_reg\[1\] _10398_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[10\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_54_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17653_ VGND VPWR VGND VPWR _10831_ keymem.prev_key1_reg\[10\] _03698_ _03670_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_72_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14865_ VPWR VGND _10330_ _10329_ keymem.prev_key0_reg\[7\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_76_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16604_ VGND VPWR VGND VPWR _02758_ _02757_ _02761_ _02759_ sky130_fd_sc_hd__a21oi_2
X_13816_ VGND VPWR VGND VPWR enc_block.block_w1_reg\[28\] _08985_ _09022_ _09286_
+ _09288_ _09287_ sky130_fd_sc_hd__a2111o_2
X_17584_ VGND VPWR VGND VPWR _02777_ _02776_ _09868_ _03644_ sky130_fd_sc_hd__a21o_2
X_14796_ _10243_ _10262_ _07386_ _10261_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_19323_ VGND VPWR _00476_ _05042_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_161_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16535_ VGND VPWR VGND VPWR _11532_ _02692_ _02694_ _11502_ sky130_fd_sc_hd__nand3_2
XFILLER_0_58_657 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13747_ VPWR VGND VGND VPWR _09091_ _09219_ _09216_ sky130_fd_sc_hd__nor2_2
XFILLER_0_39_860 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19254_ VGND VPWR _04999_ _04877_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16466_ VGND VPWR VGND VPWR _11320_ _11403_ _11204_ _11460_ _02627_ sky130_fd_sc_hd__o22a_2
X_13678_ VGND VPWR VPWR VGND _09086_ _09050_ _09071_ _09150_ sky130_fd_sc_hd__or3_2
XFILLER_0_112_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_521 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18205_ VPWR VGND _04115_ _04114_ enc_block.round_key\[108\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15417_ VPWR VGND VPWR VGND _10876_ _10877_ _10878_ _10578_ _10875_ sky130_fd_sc_hd__or4b_2
XFILLER_0_54_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12629_ VPWR VGND VPWR VGND _08184_ keymem.key_mem\[7\]\[47\] _07650_ keymem.key_mem\[9\]\[47\]
+ _07738_ _08185_ sky130_fd_sc_hd__a221o_2
X_19185_ VGND VPWR VGND VPWR _04957_ keymem.key_mem_we _03068_ _04924_ _00423_ sky130_fd_sc_hd__a31o_2
X_16397_ VGND VPWR VPWR VGND _11174_ _11338_ _11263_ _02559_ sky130_fd_sc_hd__or3_2
XFILLER_0_13_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18136_ VPWR VGND VGND VPWR _04052_ _04004_ _11057_ sky130_fd_sc_hd__nand2_2
XFILLER_0_83_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_207_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15348_ _10487_ _10810_ _10809_ _10672_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_147_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18067_ VPWR VGND VGND VPWR _03988_ _03983_ _03986_ sky130_fd_sc_hd__nand2_2
XFILLER_0_110_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_123_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15279_ VGND VPWR VPWR VGND _10286_ _10741_ key[137] _10742_ sky130_fd_sc_hd__mux2_2
XFILLER_0_257_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17018_ VGND VPWR _03142_ _02771_ _02772_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_110_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_95_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_460 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18969_ VPWR VGND VGND VPWR _04802_ _04803_ _04382_ sky130_fd_sc_hd__nor2_2
XFILLER_0_226_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_806 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_213_508 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21980_ VPWR VGND keymem.key_mem\[3\]\[54\] _06470_ _06469_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_241_828 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_94_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_154_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_187 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_256_1089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_158_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20931_ VGND VPWR VPWR VGND _01215_ _05824_ _03286_ _08922_ _05911_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_90_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1343 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23650_ keymem.prev_key0_reg\[6\] clk _00147_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20862_ VGND VPWR VPWR VGND _05867_ _04941_ keymem.key_mem\[7\]\[43\] _05875_ sky130_fd_sc_hd__mux2_2
XFILLER_0_7_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_117_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22601_ VGND VPWR _06777_ _06696_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23581_ VGND VPWR VPWR VGND clk _00082_ reset_n keymem.key_mem\[14\]\[70\] sky130_fd_sc_hd__dfrtp_2
X_20793_ VGND VPWR _01151_ _05837_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_37_819 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_92_1_Right_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25320_ VGND VPWR VPWR VGND clk _01813_ reset_n keymem.key_mem\[2\]\[33\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_8_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22532_ VGND VPWR _06754_ _06696_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_8_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_130_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1130 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25251_ VGND VPWR VPWR VGND clk _01744_ reset_n keymem.key_mem\[3\]\[92\] sky130_fd_sc_hd__dfrtp_2
X_22463_ VGND VPWR _01933_ _06725_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_165_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24202_ VGND VPWR VPWR VGND clk _00695_ reset_n keymem.key_mem\[11\]\[67\] sky130_fd_sc_hd__dfrtp_2
X_21414_ VGND VPWR VPWR VGND _06162_ _03015_ keymem.key_mem\[5\]\[46\] _06168_ sky130_fd_sc_hd__mux2_2
XFILLER_0_60_822 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22394_ VGND VPWR _01901_ _06688_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25182_ VGND VPWR VPWR VGND clk _01675_ reset_n keymem.key_mem\[3\]\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_165_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24133_ VGND VPWR VPWR VGND clk _00626_ reset_n keymem.key_mem\[12\]\[126\] sky130_fd_sc_hd__dfrtp_2
X_21345_ VGND VPWR VPWR VGND _06128_ _11039_ keymem.key_mem\[5\]\[13\] _06132_ sky130_fd_sc_hd__mux2_2
XFILLER_0_62_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_579 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_124_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24064_ VGND VPWR VPWR VGND clk _00557_ reset_n keymem.key_mem\[12\]\[57\] sky130_fd_sc_hd__dfrtp_2
X_21276_ VGND VPWR VPWR VGND _06087_ _03555_ keymem.key_mem\[6\]\[110\] _06094_ sky130_fd_sc_hd__mux2_2
X_20227_ VGND VPWR _00885_ _05537_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23015_ VGND VPWR _06976_ _06924_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_229_663 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_102_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_1188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20158_ VGND VPWR VPWR VGND _05493_ _03485_ keymem.key_mem\[10\]\[99\] _05499_ sky130_fd_sc_hd__mux2_2
XFILLER_0_244_655 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1088 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_176_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24966_ VGND VPWR VPWR VGND clk _01459_ reset_n keymem.key_mem\[5\]\[63\] sky130_fd_sc_hd__dfrtp_2
X_12980_ VPWR VGND VPWR VGND _08501_ keymem.key_mem\[14\]\[81\] _07706_ keymem.key_mem\[8\]\[81\]
+ _08265_ _08502_ sky130_fd_sc_hd__a221o_2
X_20089_ VGND VPWR VPWR VGND _05457_ _03209_ keymem.key_mem\[10\]\[66\] _05463_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_139_1_Left_406 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_243_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_188_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23917_ VGND VPWR VPWR VGND clk _00410_ reset_n keymem.key_mem\[13\]\[38\] sky130_fd_sc_hd__dfrtp_2
X_11931_ VGND VPWR _07534_ _07533_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_73_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24897_ VGND VPWR VPWR VGND clk _01390_ reset_n keymem.key_mem\[6\]\[122\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_262_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14650_ VPWR VGND VPWR VGND _10115_ _10116_ _10117_ _10113_ _10114_ sky130_fd_sc_hd__or4b_2
XFILLER_0_252_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1057 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11862_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[2\] dec_new_block\[98\]
+ _07495_ sky130_fd_sc_hd__mux2_2
X_23848_ VGND VPWR VPWR VGND clk _00341_ reset_n enc_block.block_w2_reg\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_86_229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_79_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13601_ VGND VPWR VPWR VGND _09056_ _09073_ _09071_ _09072_ _09052_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_213_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14581_ VPWR VGND VGND VPWR _09381_ _10049_ _09378_ sky130_fd_sc_hd__nor2_2
X_11793_ VGND VPWR result[63] _07460_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23779_ VGND VPWR VPWR VGND clk _00272_ reset_n enc_block.round\[3\] sky130_fd_sc_hd__dfrtp_2
X_16320_ VGND VPWR VPWR VGND _10091_ key[149] keymem.prev_key1_reg\[21\] _02483_ sky130_fd_sc_hd__mux2_2
XFILLER_0_27_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13532_ VGND VPWR VGND VPWR _09004_ _08996_ _08994_ keymem.prev_key1_reg\[4\] _09003_
+ _09002_ sky130_fd_sc_hd__a32o_2
X_25518_ VGND VPWR VPWR VGND clk _02011_ reset_n keymem.key_mem\[1\]\[103\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_113_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_137_353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16251_ VGND VPWR VGND VPWR _11282_ _11352_ _11295_ _11308_ _02415_ sky130_fd_sc_hd__o22a_2
X_25449_ VGND VPWR VPWR VGND clk _01942_ reset_n keymem.key_mem\[1\]\[34\] sky130_fd_sc_hd__dfrtp_2
X_13463_ VGND VPWR _08935_ _08934_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_10_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Left_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_183_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15202_ VGND VPWR _10665_ keymem.prev_key0_reg\[9\] _10664_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_152_334 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12414_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[27\] _07586_ keymem.key_mem\[8\]\[27\]
+ _07539_ _07990_ sky130_fd_sc_hd__a22o_2
X_16182_ VGND VPWR VGND VPWR _02347_ _11290_ _11409_ _11612_ _02346_ sky130_fd_sc_hd__a211o_2
XFILLER_0_10_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_23_524 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13394_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[122\] _08027_ _08874_ _08870_ _08875_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_183_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15133_ VPWR VGND VPWR VGND _10591_ _10596_ _10597_ _10479_ _10486_ sky130_fd_sc_hd__or4b_2
XFILLER_0_263_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12345_ VPWR VGND VPWR VGND _07926_ keymem.key_mem\[13\]\[21\] _07694_ keymem.key_mem\[2\]\[21\]
+ _07646_ _07927_ sky130_fd_sc_hd__a221o_2
XFILLER_0_49_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15064_ VGND VPWR _10528_ _10524_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19941_ VGND VPWR VPWR VGND _05246_ keymem.key_mem\[11\]\[126\] _03661_ _05383_ sky130_fd_sc_hd__mux2_2
XFILLER_0_239_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_220_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12276_ VPWR VGND VPWR VGND _07862_ keymem.key_mem\[11\]\[16\] _07861_ keymem.key_mem\[4\]\[16\]
+ _07692_ _07863_ sky130_fd_sc_hd__a221o_2
X_14015_ VGND VPWR _09487_ _09486_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19872_ VGND VPWR VPWR VGND _05339_ keymem.key_mem\[11\]\[93\] _03444_ _05347_ sky130_fd_sc_hd__mux2_2
XFILLER_0_219_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_920 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_207_302 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18823_ VPWR VGND VPWR VGND _04671_ block[39] _04576_ enc_block.block_w1_reg\[7\]
+ _04666_ _04672_ sky130_fd_sc_hd__a221o_2
XFILLER_0_120_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Left_318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_262_430 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15966_ VPWR VGND VGND VPWR _11422_ _11263_ _11266_ sky130_fd_sc_hd__nand2_2
X_18754_ VPWR VGND VGND VPWR _04609_ _04603_ _04607_ sky130_fd_sc_hd__nand2_2
XFILLER_0_65_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_222_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_222_316 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_190_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17705_ VPWR VGND VPWR VGND _02686_ _03735_ keymem.prev_key0_reg\[24\] _03730_ _00165_
+ sky130_fd_sc_hd__a22o_2
X_14917_ VGND VPWR VGND VPWR _10379_ _10375_ _10381_ _10380_ sky130_fd_sc_hd__a21oi_2
X_15897_ VGND VPWR VGND VPWR _11295_ _11352_ _11241_ _11329_ _11353_ sky130_fd_sc_hd__o22a_2
X_18685_ _04545_ _04547_ _04294_ _04546_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_172_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_850 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_187_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_76_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_203_552 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14848_ VPWR VGND VPWR VGND _10034_ _10312_ _10313_ _09602_ _09913_ sky130_fd_sc_hd__or4b_2
X_17636_ VGND VPWR _00145_ _03686_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_198_Left_465 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_81_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1084 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_231_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17567_ VGND VPWR _03302_ key[122] _03629_ _09988_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_14779_ VPWR VGND VPWR VGND _10245_ _09248_ _10244_ sky130_fd_sc_hd__or2_2
XFILLER_0_187_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_85_262 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_105_75 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19306_ VPWR VGND keymem.key_mem_we _05031_ _03485_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16518_ VGND VPWR VPWR VGND _02668_ _02669_ keymem.prev_key1_reg\[120\] _02678_ sky130_fd_sc_hd__or3_2
XFILLER_0_46_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_498 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17498_ _11535_ _03569_ _08936_ _11536_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_185_1_Left_452 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_229_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_713 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_27_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16449_ VGND VPWR VGND VPWR _11141_ _11113_ _02610_ keymem.round_ctr_reg\[0\] sky130_fd_sc_hd__a21oi_2
X_19237_ VPWR VGND keymem.key_mem\[13\]\[73\] _04988_ _04979_ VPWR VGND sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_153_2_Left_624 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_746 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_27_874 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19168_ VGND VPWR _00417_ _04946_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_147_1145 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_48_1242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18119_ VPWR VGND VPWR VGND _04036_ _04032_ _04034_ sky130_fd_sc_hd__or2_2
X_19099_ VGND VPWR VGND VPWR _04904_ keymem.key_mem_we _02340_ _04896_ _00390_ sky130_fd_sc_hd__a31o_2
XFILLER_0_170_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21130_ VGND VPWR _01308_ _06017_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_83_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_909 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21061_ VGND VPWR VPWR VGND _05972_ _10661_ keymem.key_mem\[6\]\[8\] _05981_ sky130_fd_sc_hd__mux2_2
XFILLER_0_1_495 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_239_994 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20012_ VGND VPWR _00785_ _05422_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_195_1419 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24820_ VGND VPWR VPWR VGND clk _01313_ reset_n keymem.key_mem\[6\]\[45\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_891 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_94_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24751_ VGND VPWR VPWR VGND clk _01244_ reset_n keymem.key_mem\[7\]\[104\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21963_ VGND VPWR _01698_ _06460_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_59_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23702_ keymem.prev_key0_reg\[58\] clk _00199_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_55_1246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20914_ VPWR VGND keymem.key_mem\[7\]\[67\] _05903_ _05899_ VPWR VGND sky130_fd_sc_hd__and2_2
X_24682_ VGND VPWR VPWR VGND clk _01175_ reset_n keymem.key_mem\[7\]\[35\] sky130_fd_sc_hd__dfrtp_2
X_21894_ VGND VPWR VGND VPWR _06423_ keymem.key_mem_we _11099_ _06420_ _01666_ sky130_fd_sc_hd__a31o_2
XFILLER_0_136_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23633_ VGND VPWR VPWR VGND clk _00134_ reset_n keymem.key_mem\[14\]\[122\] sky130_fd_sc_hd__dfrtp_2
X_20845_ VPWR VGND keymem.key_mem\[7\]\[35\] _05866_ _05856_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_49_454 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_232_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_85_2_Left_556 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23564_ VGND VPWR VPWR VGND clk _00065_ reset_n keymem.key_mem\[14\]\[53\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_93_1_Right_694 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20776_ VGND VPWR VGND VPWR _05828_ keymem.key_mem_we _09992_ _05821_ _01143_ sky130_fd_sc_hd__a31o_2
XFILLER_0_9_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25303_ VGND VPWR VPWR VGND clk _01796_ reset_n keymem.key_mem\[2\]\[16\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_202_Left_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_130_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22515_ VGND VPWR VPWR VGND _06739_ keymem.key_mem\[1\]\[58\] _03130_ _06745_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_863 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23495_ VPWR VGND VGND VPWR _07192_ _07356_ _04292_ sky130_fd_sc_hd__nor2_2
XFILLER_0_134_323 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25234_ VGND VPWR VPWR VGND clk _01727_ reset_n keymem.key_mem\[3\]\[75\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22446_ VGND VPWR VPWR VGND _06715_ keymem.key_mem\[1\]\[17\] _11547_ _06717_ sky130_fd_sc_hd__mux2_2
XFILLER_0_91_298 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_66_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_161_153 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_161_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_165_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25165_ VGND VPWR VPWR VGND clk _01658_ reset_n keymem.key_mem\[3\]\[6\] sky130_fd_sc_hd__dfrtp_2
X_22377_ VGND VPWR _01893_ _06679_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_66_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1231 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_27_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12130_ VPWR VGND VPWR VGND _07726_ keymem.key_mem\[5\]\[6\] _07725_ keymem.key_mem\[3\]\[6\]
+ _07690_ _07727_ sky130_fd_sc_hd__a221o_2
X_24116_ VGND VPWR VPWR VGND clk _00609_ reset_n keymem.key_mem\[12\]\[109\] sky130_fd_sc_hd__dfrtp_2
X_21328_ VGND VPWR VPWR VGND _06117_ _10193_ keymem.key_mem\[5\]\[5\] _06123_ sky130_fd_sc_hd__mux2_2
X_25096_ VGND VPWR VPWR VGND clk _01589_ reset_n keymem.key_mem\[4\]\[65\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_257_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21259_ VGND VPWR VPWR VGND _06076_ _03506_ keymem.key_mem\[6\]\[102\] _06085_ sky130_fd_sc_hd__mux2_2
X_24047_ VGND VPWR VPWR VGND clk _00540_ reset_n keymem.key_mem\[12\]\[40\] sky130_fd_sc_hd__dfrtp_2
X_12061_ VPWR VGND VPWR VGND _07660_ keymem.key_mem\[6\]\[3\] _07657_ keymem.key_mem\[8\]\[3\]
+ _07655_ _07661_ sky130_fd_sc_hd__a221o_2
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1199 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_248_279 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_211_Left_478 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_102_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15820_ VPWR VGND VGND VPWR _11275_ _11276_ _11274_ sky130_fd_sc_hd__nor2_2
XFILLER_0_205_817 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_102_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_176_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15751_ VGND VPWR VGND VPWR _11207_ _11196_ _11195_ keymem.prev_key1_reg\[20\] _09003_
+ _09002_ sky130_fd_sc_hd__a32o_2
XFILLER_0_99_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12963_ VGND VPWR enc_block.round_key\[79\] _08486_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24949_ VGND VPWR VPWR VGND clk _01442_ reset_n keymem.key_mem\[5\]\[46\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_172_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14702_ VPWR VGND VGND VPWR _09033_ _10169_ _09216_ sky130_fd_sc_hd__nor2_2
X_11914_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[28\] dec_new_block\[124\]
+ _07521_ sky130_fd_sc_hd__mux2_2
X_18470_ VPWR VGND _04354_ enc_block.block_w0_reg\[7\] enc_block.block_w0_reg\[3\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_73_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15682_ VGND VPWR VGND VPWR _10751_ _10541_ _10572_ _10619_ _10981_ _11139_ sky130_fd_sc_hd__o32a_2
XFILLER_0_38_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12894_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[73\] _07806_ keymem.key_mem\[8\]\[73\]
+ _07654_ _08424_ sky130_fd_sc_hd__a22o_2
XFILLER_0_73_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17421_ VPWR VGND VPWR VGND _03503_ _10273_ _10274_ sky130_fd_sc_hd__or2_2
X_14633_ VGND VPWR _00016_ _10100_ VPWR VGND sky130_fd_sc_hd__buf_1
X_11845_ VGND VPWR result[89] _07486_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_142_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_51_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_220_Left_487 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17352_ VPWR VGND VPWR VGND _03442_ _03438_ _03437_ key[221] _10838_ _03443_ sky130_fd_sc_hd__a221o_2
X_14564_ VGND VPWR keymem.round_ctr_reg\[0\] _10003_ _10032_ _10031_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_11776_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[23\] dec_new_block\[55\]
+ _07452_ sky130_fd_sc_hd__mux2_2
X_16303_ VPWR VGND VPWR VGND _02467_ key[20] _09795_ sky130_fd_sc_hd__or2_2
X_13515_ VPWR VGND VPWR VGND _08986_ _08985_ _08984_ _08945_ enc_block.block_w2_reg\[5\]
+ _08987_ sky130_fd_sc_hd__a221o_2
X_17283_ VPWR VGND VGND VPWR _03381_ key[214] _03077_ sky130_fd_sc_hd__nand2_2
XFILLER_0_113_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14495_ VPWR VGND VGND VPWR _09145_ _09168_ _09964_ _09129_ _09178_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_82_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19022_ _04848_ _04850_ _04103_ _04849_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_10_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16234_ VGND VPWR _02399_ keymem.prev_key0_reg\[51\] keymem.prev_key0_reg\[83\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13446_ VPWR VGND VPWR VGND _08921_ keymem.key_mem_we sky130_fd_sc_hd__inv_2
XFILLER_0_148_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16165_ VPWR VGND _11589_ _11619_ _11618_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_148_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13377_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[121\] _07812_ keymem.key_mem\[9\]\[121\]
+ _07716_ _08859_ sky130_fd_sc_hd__a22o_2
XFILLER_0_11_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_152_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_84_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15116_ VGND VPWR _10580_ _10500_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_45_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1342 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_23_387 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12328_ VPWR VGND VPWR VGND _07910_ keymem.key_mem\[13\]\[20\] _07588_ keymem.key_mem\[6\]\[20\]
+ _07908_ _07911_ sky130_fd_sc_hd__a221o_2
XFILLER_0_80_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16096_ VPWR VGND VGND VPWR _11550_ key[146] _09511_ sky130_fd_sc_hd__nand2_2
XFILLER_0_267_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15047_ VGND VPWR _10511_ _10510_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19924_ VGND VPWR _00745_ _05374_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12259_ VGND VPWR VGND VPWR _07848_ _07839_ keymem.key_mem\[11\]\[14\] _07840_ _07847_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_259_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19855_ VGND VPWR VPWR VGND _05328_ keymem.key_mem\[11\]\[85\] _03374_ _05338_ sky130_fd_sc_hd__mux2_2
XFILLER_0_120_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18806_ VPWR VGND _04656_ enc_block.block_w2_reg\[30\] enc_block.block_w3_reg\[22\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_194_1430 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19786_ VGND VPWR VPWR VGND _05292_ keymem.key_mem\[11\]\[52\] _03075_ _05302_ sky130_fd_sc_hd__mux2_2
XFILLER_0_155_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1004 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_263_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_625 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16998_ VPWR VGND VPWR VGND _03124_ keymem.prev_key1_reg\[58\] sky130_fd_sc_hd__inv_2
XFILLER_0_222_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_194_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18737_ VGND VPWR _04593_ enc_block.block_w1_reg\[7\] _04592_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15949_ VGND VPWR VGND VPWR _11402_ _11314_ _11405_ _11404_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_95_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18668_ _04530_ _04532_ _04294_ _04531_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_56_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_116_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_235_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17619_ VGND VPWR _03674_ _03673_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18599_ VGND VPWR _04470_ enc_block.block_w1_reg\[25\] _04469_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_153_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_4_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_402 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20630_ VGND VPWR _01076_ _05749_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_19_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1143 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_266_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_1176 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_131_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20561_ VGND VPWR VPWR VGND _05703_ _02873_ keymem.key_mem\[8\]\[32\] _05713_ sky130_fd_sc_hd__mux2_2
XFILLER_0_6_521 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22300_ VGND VPWR _01856_ _06639_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23280_ VPWR VGND _07164_ _07163_ enc_block.round_key\[7\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_264_1144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20492_ VGND VPWR _05676_ _05675_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_166_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_14_321 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_332 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_162_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22231_ VGND VPWR _01823_ _06603_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_48_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_836 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22162_ VPWR VGND VGND VPWR _06567_ _08933_ _05385_ sky130_fd_sc_hd__nand2_2
XFILLER_0_242_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_858 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_30_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21113_ VGND VPWR VPWR VGND _06007_ _02873_ keymem.key_mem\[6\]\[32\] _06009_ sky130_fd_sc_hd__mux2_2
XFILLER_0_242_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22093_ VGND VPWR _01759_ _06529_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_245_216 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21044_ VGND VPWR _05972_ _05971_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_103_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_201_1172 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24803_ VGND VPWR VPWR VGND clk _01296_ reset_n keymem.key_mem\[6\]\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_213_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25783_ keymem.prev_key1_reg\[99\] clk _02276_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22995_ VGND VPWR VGND VPWR _02226_ _06964_ _06954_ keymem.prev_key1_reg\[49\] sky130_fd_sc_hd__o21a_2
XFILLER_0_202_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_173_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_989 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_198_359 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24734_ VGND VPWR VPWR VGND clk _01227_ reset_n keymem.key_mem\[7\]\[87\] sky130_fd_sc_hd__dfrtp_2
X_21946_ VGND VPWR VPWR VGND _06449_ _04931_ keymem.key_mem\[3\]\[38\] _06452_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_903 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24665_ VGND VPWR VPWR VGND clk _01158_ reset_n keymem.key_mem\[7\]\[18\] sky130_fd_sc_hd__dfrtp_2
X_21877_ VGND VPWR VGND VPWR _06414_ keymem.key_mem_we _10284_ _06404_ _01658_ sky130_fd_sc_hd__a31o_2
XFILLER_0_16_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_38_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23616_ VGND VPWR VPWR VGND clk _00117_ reset_n keymem.key_mem\[14\]\[105\] sky130_fd_sc_hd__dfrtp_2
X_11630_ VPWR VGND _07369_ _07371_ _07370_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_38_947 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20828_ VPWR VGND keymem.key_mem\[7\]\[27\] _05857_ _05856_ VPWR VGND sky130_fd_sc_hd__and2_2
X_24596_ VGND VPWR VPWR VGND clk _01089_ reset_n keymem.key_mem\[8\]\[77\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_110_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_370 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23547_ VGND VPWR VPWR VGND clk _00048_ reset_n keymem.key_mem\[14\]\[36\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_94_1_Right_695 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20759_ VGND VPWR _01138_ _05816_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_52_405 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13300_ VPWR VGND VPWR VGND keymem.key_mem\[4\]\[113\] _07734_ keymem.key_mem\[1\]\[113\]
+ _07558_ _08790_ sky130_fd_sc_hd__a22o_2
XFILLER_0_110_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14280_ VGND VPWR VGND VPWR _09396_ _09411_ _09312_ _09749_ _09750_ sky130_fd_sc_hd__o22a_2
X_23478_ VGND VPWR _07341_ enc_block.round_key\[28\] _07340_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_33_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_134_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25217_ VGND VPWR VPWR VGND clk _01710_ reset_n keymem.key_mem\[3\]\[58\] sky130_fd_sc_hd__dfrtp_2
X_13231_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[106\] _07725_ keymem.key_mem\[3\]\[106\]
+ _08009_ _08728_ sky130_fd_sc_hd__a22o_2
XFILLER_0_180_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22429_ VGND VPWR _01916_ _06708_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_61_983 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_33_685 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_32_173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13162_ VPWR VGND VPWR VGND _08665_ keymem.key_mem\[14\]\[99\] _07963_ keymem.key_mem\[6\]\[99\]
+ _08137_ _08666_ sky130_fd_sc_hd__a221o_2
X_25148_ VGND VPWR VPWR VGND clk _01641_ reset_n keymem.key_mem\[4\]\[117\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12113_ VGND VPWR enc_block.round_key\[5\] _07710_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_27_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17970_ VGND VPWR _00254_ _03911_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13093_ VGND VPWR VGND VPWR _08604_ _08150_ keymem.key_mem\[3\]\[92\] _08601_ _08603_
+ sky130_fd_sc_hd__a211o_2
X_25079_ VGND VPWR VPWR VGND clk _01572_ reset_n keymem.key_mem\[4\]\[48\] sky130_fd_sc_hd__dfrtp_2
X_16921_ VPWR VGND VGND VPWR _03055_ key[178] _02875_ sky130_fd_sc_hd__nand2_2
XFILLER_0_236_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12044_ VGND VPWR _07644_ _07533_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_229_290 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19640_ VGND VPWR _00612_ _05223_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16852_ VGND VPWR _10378_ keymem.prev_key1_reg\[44\] _02992_ keymem.prev_key1_reg\[76\]
+ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_219_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15803_ VPWR VGND VPWR VGND _11173_ _11258_ _11180_ _11233_ _11259_ sky130_fd_sc_hd__or4_2
X_16783_ VGND VPWR VGND VPWR _02929_ _02928_ _02927_ key[38] sky130_fd_sc_hd__o21a_2
X_19571_ VPWR VGND keymem.key_mem\[12\]\[79\] _05188_ _05173_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13995_ VGND VPWR VGND VPWR _09389_ _09333_ _09467_ _09466_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_189_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15734_ VGND VPWR VGND VPWR enc_block.block_w2_reg\[22\] _09269_ _10387_ _11188_
+ _11190_ _11189_ sky130_fd_sc_hd__a2111o_2
X_18522_ VGND VPWR _04401_ enc_block.block_w3_reg\[8\] enc_block.block_w3_reg\[15\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_189_359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12946_ VPWR VGND VPWR VGND _08470_ keymem.key_mem\[5\]\[78\] _07725_ keymem.key_mem\[8\]\[78\]
+ _07541_ _08471_ sky130_fd_sc_hd__a221o_2
XFILLER_0_62_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_28 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15665_ VGND VPWR VGND VPWR _10609_ _10633_ _10629_ _10498_ _11122_ sky130_fd_sc_hd__o22a_2
X_18453_ VPWR VGND VGND VPWR _04328_ _04339_ _04005_ sky130_fd_sc_hd__nor2_2
X_12877_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[71\] _07597_ keymem.key_mem\[3\]\[71\]
+ _08216_ _08409_ sky130_fd_sc_hd__a22o_2
XFILLER_0_213_1043 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1065 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_200_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17404_ VGND VPWR VGND VPWR _03488_ _03221_ _02342_ _03487_ _10190_ sky130_fd_sc_hd__a211o_2
X_14616_ VGND VPWR VGND VPWR key[4] _09930_ _10083_ _10082_ _10084_ sky130_fd_sc_hd__o22a_2
X_11828_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[17\] dec_new_block\[81\]
+ _07478_ sky130_fd_sc_hd__mux2_2
X_18384_ VGND VPWR _04277_ enc_block.block_w3_reg\[5\] _04032_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15596_ VGND VPWR VPWR VGND _11053_ _11054_ _10371_ _11048_ _11049_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_44_906 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17335_ VGND VPWR VPWR VGND _03384_ keymem.key_mem\[14\]\[91\] _03427_ _03428_ sky130_fd_sc_hd__mux2_2
X_14547_ VPWR VGND VPWR VGND _09078_ _09935_ _09961_ _10014_ _10015_ sky130_fd_sc_hd__or4_2
X_11759_ VGND VPWR result[46] _07443_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17266_ VGND VPWR _00096_ _03365_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14478_ VPWR VGND VPWR VGND _09943_ _09946_ _09944_ _09942_ _09947_ sky130_fd_sc_hd__or4_2
XFILLER_0_148_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16217_ VPWR VGND VPWR VGND _11515_ _02381_ _02379_ _02378_ _02382_ sky130_fd_sc_hd__or4_2
XFILLER_0_52_950 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19005_ VGND VPWR _04835_ enc_block.round_key\[58\] _04834_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_102_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13429_ VGND VPWR VGND VPWR _07542_ keymem.key_mem\[8\]\[126\] _08903_ _08905_ _08906_
+ _07573_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_3_535 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17197_ VPWR VGND VGND VPWR _03304_ key[205] _03077_ sky130_fd_sc_hd__nand2_2
XFILLER_0_109_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1381 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16148_ VPWR VGND VPWR VGND _11601_ _11309_ _11602_ _11421_ _11528_ sky130_fd_sc_hd__or4b_2
XFILLER_0_84_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16079_ VPWR VGND VPWR VGND _11534_ keymem.prev_key0_reg\[113\] sky130_fd_sc_hd__inv_2
XFILLER_0_45_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19907_ VGND VPWR _00737_ _05365_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_209_942 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_196_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19838_ VGND VPWR _00704_ _05329_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_196_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_411 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_155_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19769_ VGND VPWR _00671_ _05293_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_159_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21800_ VGND VPWR _01624_ _06371_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_155_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22780_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[88\] _06850_ _06849_ _05013_ _02124_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_116_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21731_ VGND VPWR _01591_ _06335_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_8_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24450_ VGND VPWR VPWR VGND clk _00943_ reset_n keymem.key_mem\[9\]\[59\] sky130_fd_sc_hd__dfrtp_2
X_21662_ VGND VPWR _01558_ _06299_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23401_ VPWR VGND VGND VPWR _07192_ _07273_ _04191_ sky130_fd_sc_hd__nor2_2
X_20613_ VGND VPWR _01068_ _05740_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24381_ VGND VPWR VPWR VGND clk _00874_ reset_n keymem.key_mem\[10\]\[118\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_62_714 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21593_ VGND VPWR _06263_ _06262_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_61_202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23332_ VPWR VGND VPWR VGND _07210_ _04874_ _07209_ enc_block.block_w3_reg\[12\]
+ _07115_ _02317_ sky130_fd_sc_hd__a221o_2
X_20544_ VGND VPWR _01035_ _05704_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_166_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23263_ VPWR VGND _07148_ enc_block.block_w0_reg\[22\] enc_block.block_w3_reg\[30\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_104_326 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_171_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_148_1_Left_415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_116_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_127_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20475_ VGND VPWR VPWR VGND _05660_ _03620_ keymem.key_mem\[9\]\[120\] _05667_ sky130_fd_sc_hd__mux2_2
XFILLER_0_28_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25002_ VGND VPWR VPWR VGND clk _01495_ reset_n keymem.key_mem\[5\]\[99\] sky130_fd_sc_hd__dfrtp_2
X_22214_ VGND VPWR _01815_ _06594_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23194_ VGND VPWR _07085_ enc_block.block_w1_reg\[8\] enc_block.block_w0_reg\[16\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22145_ VGND VPWR VPWR VGND _06554_ _09991_ keymem.key_mem\[2\]\[3\] _06558_ sky130_fd_sc_hd__mux2_2
XFILLER_0_218_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_98_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22076_ VGND VPWR _01751_ _06520_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_234_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21027_ VGND VPWR VPWR VGND _05956_ _05077_ keymem.key_mem\[7\]\[121\] _05962_ sky130_fd_sc_hd__mux2_2
X_25835_ VGND VPWR VPWR VGND clk _02328_ reset_n enc_block.block_w3_reg\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_138_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_130_2_Right_202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12800_ VGND VPWR VGND VPWR _08340_ _07877_ keymem.key_mem\[10\]\[63\] _08337_ _08339_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_173_1344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13780_ VPWR VGND VPWR VGND _09252_ enc_block.block_w0_reg\[27\] _08995_ sky130_fd_sc_hd__or2_2
XFILLER_0_39_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25766_ keymem.prev_key1_reg\[82\] clk _02259_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22978_ VGND VPWR _06954_ _06881_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_230_948 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_74_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_134_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24717_ VGND VPWR VPWR VGND clk _01210_ reset_n keymem.key_mem\[7\]\[70\] sky130_fd_sc_hd__dfrtp_2
X_12731_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[56\] _08259_ _08277_ _08273_ _08278_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_201_138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21929_ VGND VPWR VGND VPWR _06442_ keymem.key_mem_we _02839_ _06432_ _01682_ sky130_fd_sc_hd__a31o_2
X_25697_ keymem.prev_key1_reg\[13\] clk _02190_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_35_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15450_ VGND VPWR VGND VPWR _10907_ _10906_ _10910_ _10911_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_32_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_338 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12662_ VGND VPWR VGND VPWR _07780_ keymem.key_mem\[5\]\[50\] _08212_ _08214_ _08215_
+ _08069_ sky130_fd_sc_hd__a2111o_2
X_24648_ VGND VPWR VPWR VGND clk _01141_ reset_n keymem.key_mem\[7\]\[1\] sky130_fd_sc_hd__dfrtp_2
X_14401_ VGND VPWR _09869_ _09866_ _09870_ _09867_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_194_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15381_ VGND VPWR VGND VPWR _10411_ _10504_ _10484_ _10566_ _10842_ sky130_fd_sc_hd__o22a_2
XFILLER_0_249_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12593_ VPWR VGND VPWR VGND _08152_ keymem.key_mem\[11\]\[43\] _08011_ keymem.key_mem\[10\]\[43\]
+ _07743_ _08153_ sky130_fd_sc_hd__a221o_2
X_24579_ VGND VPWR VPWR VGND clk _01072_ reset_n keymem.key_mem\[8\]\[60\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_25_405 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_37_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_245_Right_114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17120_ VGND VPWR _03235_ _03234_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14332_ VGND VPWR VGND VPWR _09801_ _09181_ _09059_ _09800_ _09802_ sky130_fd_sc_hd__a31o_2
XPHY_EDGE_ROW_95_1_Right_696 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_184_1440 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_184_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17051_ VGND VPWR _03173_ _03172_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14263_ VGND VPWR VGND VPWR _09563_ _09305_ _09431_ _09733_ sky130_fd_sc_hd__a21o_2
XFILLER_0_34_961 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_132_1_Left_399 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_145_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16002_ VGND VPWR VPWR VGND _11456_ _11455_ key[145] _11457_ sky130_fd_sc_hd__mux2_2
X_13214_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[104\] _08124_ _08712_ _08706_ _08713_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_81_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14194_ VPWR VGND VPWR VGND _09665_ _09189_ _09123_ sky130_fd_sc_hd__or2_2
XFILLER_0_20_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13145_ VGND VPWR enc_block.round_key\[97\] _08650_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_42_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17953_ VGND VPWR VGND VPWR _03541_ keymem.prev_key1_reg\[108\] _03900_ _10371_ sky130_fd_sc_hd__a21bo_2
X_13076_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[91\] _07918_ keymem.key_mem\[8\]\[91\]
+ _07654_ _08588_ sky130_fd_sc_hd__a22o_2
XFILLER_0_40_1131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16904_ VPWR VGND VPWR VGND _03039_ keymem.prev_key1_reg\[49\] sky130_fd_sc_hd__inv_2
X_12027_ VGND VPWR enc_block.round_key\[1\] _07628_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_194_1_Left_461 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17884_ VGND VPWR _03381_ _03852_ _03853_ _03738_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_19623_ VGND VPWR _00604_ _05214_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_206_956 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_162_2_Left_633 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16835_ VPWR VGND VPWR VGND _02976_ key[43] _08936_ sky130_fd_sc_hd__or2_2
XFILLER_0_156_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19554_ VGND VPWR VGND VPWR _05178_ keymem.key_mem_we _03252_ _05164_ _00571_ sky130_fd_sc_hd__a31o_2
XFILLER_0_156_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13978_ VGND VPWR _09450_ _09449_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_73_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16766_ VGND VPWR VPWR VGND _02884_ keymem.key_mem\[14\]\[36\] _02913_ _02914_ sky130_fd_sc_hd__mux2_2
XFILLER_0_92_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18505_ VGND VPWR _04386_ _04383_ _04385_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15717_ VGND VPWR _11173_ _11172_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12929_ VPWR VGND VPWR VGND _08455_ keymem.key_mem\[5\]\[76\] _08052_ keymem.key_mem\[8\]\[76\]
+ _08265_ _08456_ sky130_fd_sc_hd__a221o_2
XFILLER_0_232_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19485_ VGND VPWR VPWR VGND _05138_ _04933_ keymem.key_mem\[12\]\[39\] _05142_ sky130_fd_sc_hd__mux2_2
X_16697_ VGND VPWR _02850_ _02847_ _02849_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_722 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18436_ VPWR VGND VPWR VGND _04323_ _04318_ _04322_ sky130_fd_sc_hd__or2_2
XFILLER_0_237_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15648_ VPWR VGND _11105_ _11104_ keymem.prev_key1_reg\[111\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_185_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_267_1537 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_189_1362 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_7_126 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18367_ VPWR VGND VPWR VGND _04262_ _04010_ _04260_ sky130_fd_sc_hd__or2_2
X_15579_ VGND VPWR VPWR VGND _11035_ _11034_ _11038_ _10281_ _11037_ sky130_fd_sc_hd__o211a_2
XFILLER_0_111_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17318_ VPWR VGND VGND VPWR _10287_ _03412_ key[218] sky130_fd_sc_hd__nor2_2
XFILLER_0_83_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18298_ VPWR VGND _04200_ _04199_ enc_block.round_key\[116\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_17249_ VGND VPWR VGND VPWR _02396_ keymem.prev_key0_reg\[83\] _03350_ _08937_ sky130_fd_sc_hd__nand3_2
XFILLER_0_189_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_321 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_259_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_460 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20260_ VGND VPWR _00901_ _05554_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_124_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_387 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_243_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20191_ VGND VPWR _00870_ _05516_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_11_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_204_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_2_Left_565 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23950_ VGND VPWR VPWR VGND clk _00443_ reset_n keymem.key_mem\[13\]\[71\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_1355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_215_219 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_47_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22901_ VGND VPWR _02190_ _06906_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_100_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23881_ VGND VPWR VPWR VGND clk _00374_ reset_n keymem.key_mem\[13\]\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_251_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25620_ VGND VPWR VPWR VGND clk _02113_ reset_n keymem.key_mem\[0\]\[77\] sky130_fd_sc_hd__dfrtp_2
X_22832_ VGND VPWR VGND VPWR keymem.rcon_reg\[0\] _06862_ keymem.rcon_logic.tmp_rcon\[0\]
+ _06863_ _02164_ sky130_fd_sc_hd__o22a_2
XFILLER_0_195_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_56_1171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25551_ VGND VPWR VPWR VGND clk _02044_ reset_n keymem.key_mem\[0\]\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22763_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[78\] _06837_ _06836_ _04997_ _02114_
+ sky130_fd_sc_hd__a22o_2
X_24502_ VGND VPWR VPWR VGND clk _00995_ reset_n keymem.key_mem\[9\]\[111\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_52_1046 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_93_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21714_ VGND VPWR _01583_ _06326_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_220_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_211_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25482_ VGND VPWR VPWR VGND clk _01975_ reset_n keymem.key_mem\[1\]\[67\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_52_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22694_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[36\] _06790_ _06789_ _04927_ _02072_
+ sky130_fd_sc_hd__a22o_2
X_24433_ VGND VPWR VPWR VGND clk _00926_ reset_n keymem.key_mem\[9\]\[42\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_211_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21645_ VGND VPWR _01550_ _06290_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_176_395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_240_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_382 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24364_ VGND VPWR VPWR VGND clk _00857_ reset_n keymem.key_mem\[10\]\[101\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_227_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21576_ VGND VPWR _01519_ _06252_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_209_1410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_950 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23315_ VPWR VGND _07195_ enc_block.block_w1_reg\[15\] enc_block.block_w1_reg\[10\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_6_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20527_ VGND VPWR _01027_ _05695_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24295_ VGND VPWR VPWR VGND clk _00788_ reset_n keymem.key_mem\[10\]\[32\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_15_460 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_31_931 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23246_ VPWR VGND VGND VPWR _07133_ _07128_ _07132_ sky130_fd_sc_hd__nand2_2
XFILLER_0_249_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20458_ VGND VPWR VPWR VGND _05649_ _03567_ keymem.key_mem\[9\]\[112\] _05658_ sky130_fd_sc_hd__mux2_2
XFILLER_0_30_441 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_28_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23177_ VGND VPWR VPWR VGND _07054_ _07074_ keymem.prev_key1_reg\[121\] _07075_ sky130_fd_sc_hd__mux2_2
X_20389_ VGND VPWR VPWR VGND _05614_ _03322_ keymem.key_mem\[9\]\[79\] _05622_ sky130_fd_sc_hd__mux2_2
XFILLER_0_24_1137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_203_1042 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22128_ VGND VPWR _01776_ _06547_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_98_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1086 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_140_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14950_ VGND VPWR _10414_ _10413_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22059_ VGND VPWR VGND VPWR _06511_ keymem.key_mem_we _03427_ _06498_ _01743_ sky130_fd_sc_hd__a31o_2
X_13901_ VPWR VGND VGND VPWR _09373_ _09319_ _09304_ sky130_fd_sc_hd__nand2_2
X_14881_ _09044_ _10346_ _09043_ _09045_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_216_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_443 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13832_ VGND VPWR _09304_ _09261_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16620_ VGND VPWR VGND VPWR _02768_ keymem.prev_key1_reg\[124\] _02776_ _02767_ sky130_fd_sc_hd__nand3_2
X_25818_ VGND VPWR VPWR VGND clk _02311_ reset_n enc_block.block_w3_reg\[6\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_131_2_Right_203 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_138_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_806 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16551_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[121\] _02697_ _02710_ _02698_ sky130_fd_sc_hd__a21bo_2
X_13763_ VPWR VGND VGND VPWR _09149_ _09235_ _09153_ sky130_fd_sc_hd__nor2_2
XFILLER_0_69_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25749_ keymem.prev_key1_reg\[65\] clk _02242_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_35_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15502_ VGND VPWR VPWR VGND keymem.round_ctr_reg\[0\] _10961_ _10917_ _10962_ sky130_fd_sc_hd__mux2_2
X_12714_ VPWR VGND VPWR VGND _08261_ keymem.key_mem\[5\]\[55\] _07811_ keymem.key_mem\[14\]\[55\]
+ _08032_ _08262_ sky130_fd_sc_hd__a221o_2
XFILLER_0_214_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16482_ VGND VPWR VGND VPWR _02641_ _02640_ _02642_ _02643_ sky130_fd_sc_hd__a21o_2
X_19270_ VGND VPWR VPWR VGND _04993_ _05008_ keymem.key_mem\[13\]\[85\] _05009_ sky130_fd_sc_hd__mux2_2
X_13694_ VPWR VGND VPWR VGND _09044_ _09015_ _09045_ _09001_ _09166_ sky130_fd_sc_hd__or4_2
X_18221_ VGND VPWR _04129_ enc_block.block_w2_reg\[13\] _04128_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15433_ VGND VPWR VPWR VGND _10839_ _10893_ keymem.prev_key0_reg\[107\] _10894_ sky130_fd_sc_hd__or3_2
XFILLER_0_214_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_167_384 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12645_ VGND VPWR VGND VPWR _08200_ _07731_ keymem.key_mem\[13\]\[48\] _08197_ _08199_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_127_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_522 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18152_ VGND VPWR _04066_ enc_block.block_w1_reg\[16\] enc_block.block_w0_reg\[24\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_182_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15364_ VGND VPWR VGND VPWR _10826_ _09722_ _09796_ key[10] sky130_fd_sc_hd__o21a_2
XFILLER_0_65_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12576_ VGND VPWR _08137_ _07656_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_80_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_182_387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14315_ VGND VPWR VGND VPWR _09480_ _09343_ _09441_ _09349_ _09785_ sky130_fd_sc_hd__o22a_2
X_17103_ VPWR VGND VPWR VGND _03219_ key[196] sky130_fd_sc_hd__inv_2
X_18083_ VPWR VGND _04003_ _04002_ enc_block.round_key\[98\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15295_ VGND VPWR VGND VPWR _10628_ _10489_ _10609_ _10511_ _10757_ sky130_fd_sc_hd__o22a_2
XPHY_EDGE_ROW_96_1_Right_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_135_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_920 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17034_ VGND VPWR VGND VPWR _02804_ _02803_ _03157_ _03156_ sky130_fd_sc_hd__a21oi_2
X_14246_ VGND VPWR _09717_ _09516_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_1_814 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_106_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14177_ VGND VPWR VGND VPWR _09137_ _08999_ _09221_ _09080_ _09648_ sky130_fd_sc_hd__o22a_2
XFILLER_0_1_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_265_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13128_ VPWR VGND VPWR VGND _08634_ keymem.key_mem\[10\]\[96\] _07562_ keymem.key_mem\[4\]\[96\]
+ _08077_ _08635_ sky130_fd_sc_hd__a221o_2
X_18985_ VPWR VGND VPWR VGND _04817_ _04591_ _04815_ sky130_fd_sc_hd__or2_2
XFILLER_0_264_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17936_ VGND VPWR _00243_ _03888_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13059_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[89\] _08391_ keymem.key_mem\[4\]\[89\]
+ _07692_ _08573_ sky130_fd_sc_hd__a22o_2
XFILLER_0_187_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17867_ VGND VPWR _00221_ _03841_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_108_64 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_233_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19606_ VGND VPWR VPWR VGND _05205_ _05024_ keymem.key_mem\[12\]\[96\] _05206_ sky130_fd_sc_hd__mux2_2
XFILLER_0_255_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16818_ VGND VPWR VPWR VGND _09523_ key[169] keymem.prev_key1_reg\[41\] _02961_ sky130_fd_sc_hd__mux2_2
XFILLER_0_117_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17798_ VGND VPWR _03795_ _03794_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19537_ VGND VPWR VGND VPWR _05169_ keymem.key_mem_we _03184_ _05164_ _00563_ sky130_fd_sc_hd__a31o_2
XFILLER_0_191_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16749_ VGND VPWR VPWR VGND _09928_ _02897_ _02896_ _02898_ sky130_fd_sc_hd__mux2_2
XFILLER_0_117_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_191_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_75_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19468_ VGND VPWR VGND VPWR _05132_ keymem.key_mem_we _02862_ _05121_ _00531_ sky130_fd_sc_hd__a31o_2
XFILLER_0_18_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1282 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_57_850 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_947 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_124_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_552 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18419_ VGND VPWR _04307_ enc_block.block_w1_reg\[31\] enc_block.block_w0_reg\[7\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19399_ VGND VPWR _05095_ _05094_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_29_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_267_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_382 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21430_ VGND VPWR _01449_ _06176_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_12_1085 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21361_ VGND VPWR _06140_ _06116_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_31_216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_226_1031 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23100_ VGND VPWR VPWR VGND _06992_ _07026_ keymem.prev_key1_reg\[92\] _07027_ sky130_fd_sc_hd__mux2_2
XFILLER_0_140_95 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20312_ VGND VPWR VPWR VGND _05580_ _02972_ keymem.key_mem\[9\]\[42\] _05582_ sky130_fd_sc_hd__mux2_2
XFILLER_0_47_1159 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_128_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24080_ VGND VPWR VPWR VGND clk _00573_ reset_n keymem.key_mem\[12\]\[73\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_226_1064 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21292_ VGND VPWR _01385_ _06102_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_25_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23031_ VGND VPWR VGND VPWR _06985_ _03199_ _03198_ _03201_ _06951_ sky130_fd_sc_hd__a211o_2
XFILLER_0_40_772 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20243_ VGND VPWR _00893_ _05545_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_99_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20174_ VGND VPWR _00862_ _05507_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_200_1226 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_99_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_889 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_239_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24982_ VGND VPWR VPWR VGND clk _01475_ reset_n keymem.key_mem\[5\]\[79\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_1200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23933_ VGND VPWR VPWR VGND clk _00426_ reset_n keymem.key_mem\[13\]\[54\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_239_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_157_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23864_ VGND VPWR VPWR VGND clk _00357_ reset_n enc_block.block_w2_reg\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_1108 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_93_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25603_ VGND VPWR VPWR VGND clk _02096_ reset_n keymem.key_mem\[0\]\[60\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_168_115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22815_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[114\] _06860_ _06859_ _05062_ _02150_
+ sky130_fd_sc_hd__a22o_2
X_23795_ VGND VPWR VPWR VGND clk _00288_ reset_n enc_block.block_w0_reg\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_36_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25534_ VGND VPWR VPWR VGND clk _02027_ reset_n keymem.key_mem\[1\]\[119\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_211_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_66_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22746_ VGND VPWR _02103_ _06838_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_251_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_850 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_149_384 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25465_ VGND VPWR VPWR VGND clk _01958_ reset_n keymem.key_mem\[1\]\[50\] sky130_fd_sc_hd__dfrtp_2
X_22677_ VGND VPWR _02062_ _06810_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_35_500 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_47_371 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12430_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[29\] _07703_ keymem.key_mem\[14\]\[29\]
+ _08003_ _08004_ sky130_fd_sc_hd__a22o_2
X_24416_ VGND VPWR VPWR VGND clk _00909_ reset_n keymem.key_mem\[9\]\[25\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_47_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21628_ VGND VPWR _01542_ _06281_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_191_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25396_ VGND VPWR VPWR VGND clk _01889_ reset_n keymem.key_mem\[2\]\[109\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_191_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_246_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_117_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24347_ VGND VPWR VPWR VGND clk _00840_ reset_n keymem.key_mem\[10\]\[84\] sky130_fd_sc_hd__dfrtp_2
X_12361_ VGND VPWR VGND VPWR _07942_ _07629_ keymem.key_mem\[10\]\[22\] _07939_ _07941_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_63_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21559_ VGND VPWR VPWR VGND _06242_ _03585_ keymem.key_mem\[5\]\[115\] _06244_ sky130_fd_sc_hd__mux2_2
X_14100_ VGND VPWR VGND VPWR _09328_ _09571_ _09339_ _09306_ _09486_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_50_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_107_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_240 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15080_ VPWR VGND VPWR VGND _10456_ _10445_ _10444_ _10443_ _10544_ sky130_fd_sc_hd__or4_2
XFILLER_0_146_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12292_ VGND VPWR _07878_ _07752_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24278_ VGND VPWR VPWR VGND clk _00771_ reset_n keymem.key_mem\[10\]\[15\] sky130_fd_sc_hd__dfrtp_2
X_14031_ VPWR VGND VPWR VGND _09501_ _09502_ _09503_ _09498_ _09499_ sky130_fd_sc_hd__or4b_2
XFILLER_0_107_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23229_ VGND VPWR _07117_ enc_block.block_w3_reg\[26\] _07116_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_311 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_246_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18770_ VPWR VGND VPWR VGND _04623_ _04550_ _04622_ enc_block.block_w2_reg\[2\] _04602_
+ _00342_ sky130_fd_sc_hd__a221o_2
XFILLER_0_257_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15982_ VGND VPWR VGND VPWR _11383_ _11437_ _11438_ _11364_ _11406_ sky130_fd_sc_hd__nor4_2
XFILLER_0_140_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_262_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17721_ VGND VPWR VGND VPWR _03737_ keymem.prev_key1_reg\[29\] _03747_ _03738_ sky130_fd_sc_hd__a21oi_2
X_14933_ VGND VPWR VGND VPWR _10397_ _10396_ _10395_ keymem.prev_key1_reg\[8\] _08955_
+ _08942_ sky130_fd_sc_hd__a32o_2
XFILLER_0_257_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17652_ VGND VPWR _00150_ _03697_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14864_ VPWR VGND _10329_ keymem.prev_key0_reg\[71\] keymem.prev_key0_reg\[39\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_251_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_192_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_203_756 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16603_ _02758_ _02760_ _02757_ _02759_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_13815_ enc_block.sword_ctr_reg\[1\] _09287_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[28\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_14795_ VPWR VGND VGND VPWR _09438_ _10245_ _10248_ _10260_ _10261_ sky130_fd_sc_hd__and4b_2
XFILLER_0_114_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_2_Right_204 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17583_ VGND VPWR VGND VPWR _03643_ _03302_ _08937_ key[124] sky130_fd_sc_hd__o21a_2
XFILLER_0_97_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19322_ VGND VPWR VPWR VGND _05025_ _05041_ keymem.key_mem\[13\]\[104\] _05042_ sky130_fd_sc_hd__mux2_2
X_13746_ VPWR VGND VGND VPWR _09216_ _09217_ _09218_ _09089_ _09200_ sky130_fd_sc_hd__o22ai_2
X_16534_ VGND VPWR VGND VPWR _11532_ _11502_ _02692_ _02693_ sky130_fd_sc_hd__a21o_2
XFILLER_0_70_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19253_ VGND VPWR _00450_ _04998_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_151_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16465_ VGND VPWR VGND VPWR _11218_ _11318_ _11314_ _11327_ _02626_ sky130_fd_sc_hd__o22a_2
X_13677_ VGND VPWR _09149_ _09148_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_72_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18204_ VPWR VGND VPWR VGND _04113_ block[108] _04076_ enc_block.block_w2_reg\[12\]
+ _04007_ _04114_ sky130_fd_sc_hd__a221o_2
XFILLER_0_112_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15416_ VGND VPWR VGND VPWR _10521_ _10546_ _10476_ _10557_ _10877_ sky130_fd_sc_hd__o22a_2
X_12628_ VPWR VGND VPWR VGND keymem.key_mem\[8\]\[47\] _07654_ keymem.key_mem\[1\]\[47\]
+ _07624_ _08184_ sky130_fd_sc_hd__a22o_2
X_16396_ VGND VPWR VGND VPWR _11253_ _11314_ _11270_ _11345_ _02558_ sky130_fd_sc_hd__o22a_2
XFILLER_0_26_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19184_ VPWR VGND keymem.key_mem\[13\]\[51\] _04957_ _04915_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_170_302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15347_ VPWR VGND VGND VPWR _10464_ _10809_ _10463_ sky130_fd_sc_hd__nor2_2
X_18135_ VPWR VGND _04051_ _04050_ enc_block.round_key\[102\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_12559_ VPWR VGND VPWR VGND _08121_ keymem.key_mem\[14\]\[40\] _07721_ keymem.key_mem\[6\]\[40\]
+ _07712_ _08122_ sky130_fd_sc_hd__a221o_2
XFILLER_0_186_1398 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1061 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_262_1231 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_102_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18066_ VPWR VGND VPWR VGND _03987_ _03983_ _03986_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_97_1_Right_698 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15278_ VPWR VGND _10741_ keymem.prev_key1_reg\[41\] keymem.prev_key1_reg\[9\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_13_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_83_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Right_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14229_ VGND VPWR VPWR VGND _09011_ _09185_ _09089_ _09700_ sky130_fd_sc_hd__or3_2
XFILLER_0_257_417 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17017_ VGND VPWR _00071_ _03141_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_186_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_201_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_688 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_956 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18968_ VGND VPWR _04802_ _04800_ _04801_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17919_ VGND VPWR VPWR VGND _03876_ key[225] keymem.prev_key1_reg\[97\] _03877_ sky130_fd_sc_hd__mux2_2
XFILLER_0_20_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18899_ VPWR VGND VPWR VGND block[47] _03979_ enc_block.block_w0_reg\[15\] _03977_
+ _04740_ sky130_fd_sc_hd__a22o_2
X_20930_ VPWR VGND VGND VPWR _05911_ keymem.key_mem\[7\]\[75\] _05824_ sky130_fd_sc_hd__nand2_2
XFILLER_0_90_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_157_1_Left_424 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_94_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_135_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_234_1366 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20861_ VGND VPWR _01182_ _05874_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_230_1208 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22600_ VGND VPWR _06776_ _03859_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_18_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23580_ VGND VPWR VPWR VGND clk _00081_ reset_n keymem.key_mem\[14\]\[69\] sky130_fd_sc_hd__dfrtp_2
X_20792_ VGND VPWR VPWR VGND _05820_ _04894_ keymem.key_mem\[7\]\[11\] _05837_ sky130_fd_sc_hd__mux2_2
XFILLER_0_64_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22531_ VGND VPWR _06753_ _03859_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_158_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_130_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25250_ VGND VPWR VPWR VGND clk _01743_ reset_n keymem.key_mem\[3\]\[91\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_267_1142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_146_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_63_138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22462_ VGND VPWR VPWR VGND _06715_ keymem.key_mem\[1\]\[25\] _02721_ _06725_ sky130_fd_sc_hd__mux2_2
XFILLER_0_161_302 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24201_ VGND VPWR VPWR VGND clk _00694_ reset_n keymem.key_mem\[11\]\[66\] sky130_fd_sc_hd__dfrtp_2
X_21413_ VGND VPWR _01441_ _06167_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_32_503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25181_ VGND VPWR VPWR VGND clk _01674_ reset_n keymem.key_mem\[3\]\[22\] sky130_fd_sc_hd__dfrtp_2
X_22393_ VGND VPWR VPWR VGND _06680_ _03627_ keymem.key_mem\[2\]\[121\] _06688_ sky130_fd_sc_hd__mux2_2
XFILLER_0_71_182 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24132_ VGND VPWR VPWR VGND clk _00625_ reset_n keymem.key_mem\[12\]\[125\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_71_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21344_ VGND VPWR _01408_ _06131_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_249_918 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24063_ VGND VPWR VPWR VGND clk _00556_ reset_n keymem.key_mem\[12\]\[56\] sky130_fd_sc_hd__dfrtp_2
X_21275_ VGND VPWR _01377_ _06093_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_124_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23014_ VGND VPWR VPWR VGND _02234_ _03113_ _03117_ _06925_ _06975_ sky130_fd_sc_hd__o31a_2
X_20226_ VGND VPWR VPWR VGND _05535_ _09725_ keymem.key_mem\[9\]\[1\] _05537_ sky130_fd_sc_hd__mux2_2
XFILLER_0_99_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_204_1181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_141_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_243_100 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20157_ VGND VPWR _00854_ _05498_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_244_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_176_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_102_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_244_667 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24965_ VGND VPWR VPWR VGND clk _01458_ reset_n keymem.key_mem\[5\]\[62\] sky130_fd_sc_hd__dfrtp_2
X_20088_ VGND VPWR _00821_ _05462_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_89_1_Left_356 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11930_ VGND VPWR VGND VPWR _07527_ _07530_ _07532_ _07531_ _07533_ sky130_fd_sc_hd__o22a_2
X_23916_ VGND VPWR VPWR VGND clk _00409_ reset_n keymem.key_mem\[13\]\[37\] sky130_fd_sc_hd__dfrtp_2
X_24896_ VGND VPWR VPWR VGND clk _01389_ reset_n keymem.key_mem\[6\]\[121\] sky130_fd_sc_hd__dfrtp_2
X_11861_ VGND VPWR result[97] _07494_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23847_ VGND VPWR VPWR VGND clk _00340_ reset_n enc_block.block_w2_reg\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_252_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_196_243 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13600_ VPWR VGND VPWR VGND _09010_ _09039_ _08971_ _09009_ _09072_ sky130_fd_sc_hd__or4_2
XFILLER_0_39_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14580_ VPWR VGND VGND VPWR _09481_ _10047_ _09331_ _09363_ _09553_ _10048_ sky130_fd_sc_hd__a311o_2
XFILLER_0_79_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11792_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[31\] dec_new_block\[63\]
+ _07460_ sky130_fd_sc_hd__mux2_2
X_23778_ VGND VPWR VPWR VGND clk _00271_ reset_n enc_block.round\[2\] sky130_fd_sc_hd__dfrtp_2
X_13531_ VGND VPWR _09003_ _08954_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_55_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22729_ VGND VPWR _02095_ _06829_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25517_ VGND VPWR VPWR VGND clk _02010_ reset_n keymem.key_mem\[1\]\[102\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_149_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_274 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16250_ VGND VPWR VGND VPWR _11252_ _11270_ _11257_ _11465_ _02414_ sky130_fd_sc_hd__o22a_2
X_25448_ VGND VPWR VPWR VGND clk _01941_ reset_n keymem.key_mem\[1\]\[33\] sky130_fd_sc_hd__dfrtp_2
X_13462_ VPWR VGND VPWR VGND _08933_ _08934_ _07386_ keymem.round_ctr_reg\[1\] sky130_fd_sc_hd__or3b_2
XFILLER_0_137_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15201_ VGND VPWR _10664_ keymem.prev_key0_reg\[41\] keymem.prev_key0_reg\[73\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
X_12413_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[27\] _07609_ keymem.key_mem\[9\]\[27\]
+ _07738_ _07989_ sky130_fd_sc_hd__a22o_2
X_16181_ VGND VPWR VGND VPWR _11349_ _11339_ _11527_ _11283_ _02346_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_183_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25379_ VGND VPWR VPWR VGND clk _01872_ reset_n keymem.key_mem\[2\]\[92\] sky130_fd_sc_hd__dfrtp_2
X_13393_ VGND VPWR VGND VPWR _08874_ _07808_ keymem.key_mem\[12\]\[122\] _08871_ _08873_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_152_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15132_ VGND VPWR VGND VPWR _10437_ _10411_ _10595_ _10593_ _10596_ sky130_fd_sc_hd__o22a_2
XPHY_EDGE_ROW_171_2_Left_642 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12344_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[21\] _07560_ keymem.key_mem\[12\]\[21\]
+ _07577_ _07926_ sky130_fd_sc_hd__a22o_2
XFILLER_0_62_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_107_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15063_ VGND VPWR _10527_ _10526_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_49_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19940_ VGND VPWR _00753_ _05382_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12275_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[16\] _07567_ keymem.key_mem\[1\]\[16\]
+ _07556_ _07862_ sky130_fd_sc_hd__a22o_2
XFILLER_0_50_399 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14014_ VGND VPWR _09486_ _09485_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19871_ VGND VPWR _00720_ _05346_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_247_461 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18822_ VPWR VGND VGND VPWR _04670_ _04671_ _04478_ sky130_fd_sc_hd__nor2_2
XFILLER_0_219_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18753_ VPWR VGND VPWR VGND _04608_ _04603_ _04607_ sky130_fd_sc_hd__or2_2
XFILLER_0_223_807 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_179_1191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15965_ VGND VPWR VGND VPWR _11420_ _11367_ _11421_ _11204_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_257_1366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_486 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17704_ VPWR VGND VGND VPWR _03734_ _03735_ _03731_ sky130_fd_sc_hd__nor2_2
X_14916_ VGND VPWR VPWR VGND _09730_ _10372_ key[136] _10380_ sky130_fd_sc_hd__mux2_2
X_18684_ VPWR VGND VPWR VGND _04546_ _04319_ _04544_ sky130_fd_sc_hd__or2_2
X_15896_ VGND VPWR _11352_ _11351_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_118_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17635_ VGND VPWR VPWR VGND _03681_ _03685_ keymem.prev_key0_reg\[4\] _03686_ sky130_fd_sc_hd__mux2_2
X_14847_ VGND VPWR VGND VPWR _09441_ _09397_ _09431_ _09371_ _09437_ _10312_ sky130_fd_sc_hd__o32a_2
XFILLER_0_231_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_81_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_133_2_Right_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17566_ VGND VPWR _00133_ _03628_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_19_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14778_ VGND VPWR VGND VPWR _09268_ _09456_ _09475_ _09420_ _09309_ _10244_ sky130_fd_sc_hd__o32a_2
XFILLER_0_14_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19305_ VGND VPWR _00470_ _05030_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_128_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16517_ VGND VPWR _02677_ _09722_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13729_ VGND VPWR VGND VPWR _09200_ _09184_ _09201_ _09185_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_105_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17497_ VGND VPWR _00124_ _03568_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19236_ VGND VPWR _00444_ _04987_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16448_ VGND VPWR _00034_ _02609_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_27_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_886 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_229_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19167_ VGND VPWR VPWR VGND _04928_ _04945_ keymem.key_mem\[13\]\[45\] _04946_ sky130_fd_sc_hd__mux2_2
XFILLER_0_27_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16379_ VGND VPWR VGND VPWR _02541_ _02542_ _02540_ _02539_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_121_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_186_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_121_64 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18118_ VPWR VGND VGND VPWR _04035_ _04032_ _04034_ sky130_fd_sc_hd__nand2_2
XFILLER_0_48_1254 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_83_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_223_1001 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19098_ VPWR VGND keymem.key_mem\[13\]\[18\] _04904_ _04903_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_44_1118 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_83_1167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18049_ VPWR VGND VGND VPWR _09239_ _03971_ _03970_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_98_1_Right_699 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_731 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21060_ VGND VPWR _01275_ _05980_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20011_ VGND VPWR VPWR VGND _05413_ _02812_ keymem.key_mem\[10\]\[29\] _05422_ sky130_fd_sc_hd__mux2_2
XFILLER_0_39_82 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_667 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24750_ VGND VPWR VPWR VGND clk _01243_ reset_n keymem.key_mem\[7\]\[103\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_207_881 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_158_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_146_61 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21962_ VGND VPWR VPWR VGND _06449_ _04947_ keymem.key_mem\[3\]\[46\] _06460_ sky130_fd_sc_hd__mux2_2
XFILLER_0_94_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23701_ keymem.prev_key0_reg\[57\] clk _00198_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20913_ VGND VPWR _01206_ _05902_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24681_ VGND VPWR VPWR VGND clk _01174_ reset_n keymem.key_mem\[7\]\[34\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_7_1001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21893_ VPWR VGND keymem.key_mem\[3\]\[14\] _06423_ _06413_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_55_1258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23632_ VGND VPWR VPWR VGND clk _00133_ reset_n keymem.key_mem\[14\]\[121\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_7_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20844_ VGND VPWR VGND VPWR _05865_ keymem.key_mem_we _02894_ _05864_ _01174_ sky130_fd_sc_hd__a31o_2
XFILLER_0_76_230 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_7_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23563_ VGND VPWR VPWR VGND clk _00064_ reset_n keymem.key_mem\[14\]\[52\] sky130_fd_sc_hd__dfrtp_2
X_20775_ VPWR VGND keymem.key_mem\[7\]\[3\] _05828_ _05824_ VPWR VGND sky130_fd_sc_hd__and2_2
X_25302_ VGND VPWR VPWR VGND clk _01795_ reset_n keymem.key_mem\[2\]\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_18_831 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_76_296 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22514_ VGND VPWR _01965_ _06744_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_247_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23494_ VGND VPWR _07355_ enc_block.round_key\[30\] _07354_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_130_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_335 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25233_ VGND VPWR VPWR VGND clk _01726_ reset_n keymem.key_mem\[3\]\[74\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_51_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22445_ VGND VPWR _01924_ _06716_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_134_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25164_ VGND VPWR VPWR VGND clk _01657_ reset_n keymem.key_mem\[3\]\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_867 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22376_ VGND VPWR VPWR VGND _06669_ _03573_ keymem.key_mem\[2\]\[113\] _06679_ sky130_fd_sc_hd__mux2_2
XFILLER_0_165_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24115_ VGND VPWR VPWR VGND clk _00608_ reset_n keymem.key_mem\[12\]\[108\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_62_1218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_66_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21327_ VGND VPWR _01400_ _06122_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_60_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25095_ VGND VPWR VPWR VGND clk _01588_ reset_n keymem.key_mem\[4\]\[64\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_243 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24046_ VGND VPWR VPWR VGND clk _00539_ reset_n keymem.key_mem\[12\]\[39\] sky130_fd_sc_hd__dfrtp_2
X_12060_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[3\] _07659_ keymem.key_mem\[11\]\[3\]
+ _07658_ _07660_ sky130_fd_sc_hd__a22o_2
XFILLER_0_257_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21258_ VGND VPWR _01369_ _06084_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_187_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20209_ VGND VPWR _00879_ _05525_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21189_ VGND VPWR _06048_ _03227_ _01336_ _05985_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_102_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_913 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15750_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[22\] _08955_ _11206_ _08942_ _11190_
+ _11191_ sky130_fd_sc_hd__a32oi_2
X_12962_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[79\] _08449_ _08485_ _08481_ _08486_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_176_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24948_ VGND VPWR VPWR VGND clk _01441_ reset_n keymem.key_mem\[5\]\[45\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_172_1217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_73_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_172_1239 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_137_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11913_ VGND VPWR result[123] _07520_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14701_ VGND VPWR VGND VPWR _10156_ _10168_ _10166_ _10167_ _10162_ sky130_fd_sc_hd__and4bb_2
X_15681_ VGND VPWR VPWR VGND _11136_ _10514_ _11138_ _11076_ _11137_ sky130_fd_sc_hd__o211a_2
XFILLER_0_59_219 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_73_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12893_ VPWR VGND VPWR VGND _08422_ keymem.key_mem\[3\]\[73\] _07691_ keymem.key_mem\[10\]\[73\]
+ _07786_ _08423_ sky130_fd_sc_hd__a221o_2
XFILLER_0_231_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24879_ VGND VPWR VPWR VGND clk _01372_ reset_n keymem.key_mem\[6\]\[104\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_34_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_212_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17420_ VGND VPWR VPWR VGND _03029_ _03501_ key[102] _03502_ sky130_fd_sc_hd__mux2_2
X_11844_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[25\] dec_new_block\[89\]
+ _07486_ sky130_fd_sc_hd__mux2_2
X_14632_ VGND VPWR VPWR VGND _09864_ keymem.key_mem\[14\]\[4\] _10099_ _10100_ sky130_fd_sc_hd__mux2_2
XFILLER_0_206_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_169_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_28_606 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_224 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14563_ VPWR VGND VPWR VGND _10018_ _10030_ _10027_ _10012_ _10031_ sky130_fd_sc_hd__or4_2
X_17351_ VGND VPWR VPWR VGND _03440_ _03439_ _03442_ _09722_ _03441_ sky130_fd_sc_hd__o211a_2
X_11775_ VGND VPWR result[54] _07451_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_27_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_628 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_937 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16302_ VGND VPWR VGND VPWR _02464_ _02463_ _02466_ keymem.prev_key0_reg\[20\] sky130_fd_sc_hd__a21oi_2
X_13514_ enc_block.sword_ctr_reg\[1\] _08986_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[5\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_14494_ VPWR VGND VGND VPWR _09216_ _09113_ _09963_ _09156_ _09116_ sky130_fd_sc_hd__o22ai_2
X_17282_ VGND VPWR VPWR VGND _02599_ _02600_ _09868_ _03380_ sky130_fd_sc_hd__or3_2
X_19021_ VPWR VGND VPWR VGND _04849_ _04637_ _04847_ sky130_fd_sc_hd__or2_2
XFILLER_0_187_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16233_ VPWR VGND VPWR VGND _02398_ _09932_ _02396_ sky130_fd_sc_hd__or2_2
X_13445_ VGND VPWR enc_block.round_key\[127\] _08920_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_10_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_694 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_246_1056 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16164_ VPWR VGND VGND VPWR _11594_ _11608_ _11617_ _11618_ sky130_fd_sc_hd__nor3_2
XFILLER_0_84_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13376_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[121\] _07650_ keymem.key_mem\[2\]\[121\]
+ _08116_ _08858_ sky130_fd_sc_hd__a22o_2
XFILLER_0_144_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_344 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_148_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15115_ VPWR VGND VGND VPWR _10536_ _10579_ _10482_ sky130_fd_sc_hd__nor2_2
X_12327_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[20\] _07650_ keymem.key_mem\[10\]\[20\]
+ _07909_ _07910_ sky130_fd_sc_hd__a22o_2
XFILLER_0_84_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16095_ VGND VPWR _11549_ keymem.prev_key1_reg\[18\] keymem.prev_key1_reg\[50\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_146_1190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15046_ VGND VPWR _10510_ _10509_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19923_ VGND VPWR VPWR VGND _05372_ keymem.key_mem\[11\]\[117\] _03600_ _05374_ sky130_fd_sc_hd__mux2_2
XFILLER_0_43_1140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12258_ VPWR VGND VPWR VGND _07846_ keymem.key_mem\[9\]\[14\] _07842_ keymem.key_mem\[4\]\[14\]
+ _07841_ _07847_ sky130_fd_sc_hd__a221o_2
XFILLER_0_267_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19854_ VGND VPWR _00712_ _05337_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12189_ VGND VPWR _07782_ _07744_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_236_954 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_207_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18805_ VPWR VGND VPWR VGND _04655_ _04550_ _04653_ enc_block.block_w2_reg\[5\] _04602_
+ _00345_ sky130_fd_sc_hd__a221o_2
XFILLER_0_120_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_442 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19785_ VGND VPWR _00679_ _05301_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_208_689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_194_1442 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16997_ VGND VPWR VPWR VGND _03121_ _02691_ _03123_ _09514_ _03122_ sky130_fd_sc_hd__o211a_2
XFILLER_0_155_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18736_ VPWR VGND _04592_ enc_block.block_w2_reg\[24\] enc_block.block_w3_reg\[16\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_267_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15948_ VGND VPWR _11404_ _11403_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_194_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_155_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18667_ VPWR VGND VGND VPWR _04531_ _04461_ _04529_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_259_Right_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15879_ VPWR VGND VGND VPWR _11252_ _11282_ _11335_ _11334_ _11318_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_91_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_52_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_489 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17618_ VPWR VGND VGND VPWR _09637_ _02947_ _03672_ _03673_ sky130_fd_sc_hd__nor3_2
XFILLER_0_263_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18598_ VPWR VGND _04469_ enc_block.block_w2_reg\[23\] enc_block.block_w2_reg\[16\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_114_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_4_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_2_Right_206 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17549_ VGND VPWR VPWR VGND _03593_ keymem.key_mem\[14\]\[119\] _03613_ _03614_ sky130_fd_sc_hd__mux2_2
X_20560_ VGND VPWR _01043_ _05712_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_188_1279 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_27_661 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19219_ VPWR VGND keymem.key_mem_we _04977_ _03209_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_190_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20491_ VPWR VGND VGND VPWR _08921_ _05675_ _05240_ _08925_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_166_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22230_ VGND VPWR VPWR VGND _06600_ _02985_ keymem.key_mem\[2\]\[43\] _06603_ sky130_fd_sc_hd__mux2_2
XFILLER_0_162_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_1073 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_74_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22161_ VGND VPWR _01790_ _06566_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_63_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21112_ VGND VPWR _01299_ _06008_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22092_ VGND VPWR VPWR VGND _06527_ _05048_ keymem.key_mem\[3\]\[107\] _06529_ sky130_fd_sc_hd__mux2_2
XFILLER_0_1_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21043_ VGND VPWR _05971_ _05970_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_10_594 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_103_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24802_ VGND VPWR VPWR VGND clk _01295_ reset_n keymem.key_mem\[6\]\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_173_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22994_ VGND VPWR VGND VPWR _06964_ _03038_ _03037_ _03045_ _06951_ sky130_fd_sc_hd__a211o_2
X_25782_ keymem.prev_key1_reg\[98\] clk _02275_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_241_434 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_55_1000 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_173_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21945_ VGND VPWR VGND VPWR _06451_ keymem.key_mem_we _02924_ _06446_ _01689_ sky130_fd_sc_hd__a31o_2
X_24733_ VGND VPWR VPWR VGND clk _01226_ reset_n keymem.key_mem\[7\]\[86\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_253_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_213_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_692 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24664_ VGND VPWR VPWR VGND clk _01157_ reset_n keymem.key_mem\[7\]\[17\] sky130_fd_sc_hd__dfrtp_2
X_21876_ VPWR VGND keymem.key_mem\[3\]\[6\] _06414_ _06413_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_166_224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23615_ VGND VPWR VPWR VGND clk _00116_ reset_n keymem.key_mem\[14\]\[104\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20827_ VGND VPWR _05856_ _05823_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24595_ VGND VPWR VPWR VGND clk _01088_ reset_n keymem.key_mem\[8\]\[76\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_296 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23546_ VGND VPWR VPWR VGND clk _00047_ reset_n keymem.key_mem\[14\]\[35\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_64_244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20758_ VGND VPWR VPWR VGND _05679_ _03661_ keymem.key_mem\[8\]\[126\] _05816_ sky130_fd_sc_hd__mux2_2
XFILLER_0_110_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_382 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_181_238 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23477_ VPWR VGND VPWR VGND _07339_ block[28] _04139_ enc_block.block_w3_reg\[28\]
+ _04138_ _07340_ sky130_fd_sc_hd__a221o_2
X_20689_ VGND VPWR VPWR VGND _05772_ _03443_ keymem.key_mem\[8\]\[93\] _05780_ sky130_fd_sc_hd__mux2_2
X_25216_ VGND VPWR VPWR VGND clk _01709_ reset_n keymem.key_mem\[3\]\[57\] sky130_fd_sc_hd__dfrtp_2
X_13230_ VGND VPWR VGND VPWR _07835_ keymem.key_mem\[13\]\[106\] _08724_ _08726_ _08727_
+ _08599_ sky130_fd_sc_hd__a2111o_2
X_22428_ VGND VPWR VPWR VGND _06702_ keymem.key_mem\[1\]\[8\] _10662_ _06708_ sky130_fd_sc_hd__mux2_2
XFILLER_0_33_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_187 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_180_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13161_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[99\] _07612_ keymem.key_mem\[12\]\[99\]
+ _07787_ _08665_ sky130_fd_sc_hd__a22o_2
X_25147_ VGND VPWR VPWR VGND clk _01640_ reset_n keymem.key_mem\[4\]\[116\] sky130_fd_sc_hd__dfrtp_2
X_22359_ VGND VPWR _01884_ _06670_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_221_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_182_1390 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_260_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12112_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[5\] _07645_ _07709_ _07701_ _07710_
+ sky130_fd_sc_hd__o22a_2
X_13092_ VPWR VGND VPWR VGND _08602_ keymem.key_mem\[9\]\[92\] _07672_ keymem.key_mem\[4\]\[92\]
+ _07854_ _08603_ sky130_fd_sc_hd__a221o_2
X_25078_ VGND VPWR VPWR VGND clk _01571_ reset_n keymem.key_mem\[4\]\[47\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_221_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16920_ VGND VPWR VGND VPWR _03054_ _03053_ _03052_ _03051_ _09534_ sky130_fd_sc_hd__o211ai_2
X_24029_ VGND VPWR VPWR VGND clk _00522_ reset_n keymem.key_mem\[12\]\[22\] sky130_fd_sc_hd__dfrtp_2
X_12043_ VGND VPWR enc_block.round_key\[2\] _07643_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16851_ VGND VPWR VGND VPWR _10190_ _09796_ _02988_ _10963_ _02991_ sky130_fd_sc_hd__a31o_2
X_15802_ VGND VPWR _11258_ _11248_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_219_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19570_ VGND VPWR _05187_ _05092_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16782_ VGND VPWR _02928_ _09512_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13994_ VGND VPWR _09466_ _09366_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18521_ VPWR VGND _04400_ _04318_ enc_block.block_w0_reg\[1\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_137_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15733_ VGND VPWR VGND VPWR _11189_ enc_block.sword_ctr_reg\[0\] enc_block.block_w1_reg\[22\]
+ enc_block.sword_ctr_reg\[1\] sky130_fd_sc_hd__and3b_2
XFILLER_0_232_467 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_220_607 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12945_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[78\] _07618_ keymem.key_mem\[1\]\[78\]
+ _07557_ _08470_ sky130_fd_sc_hd__a22o_2
X_18452_ VPWR VGND _04338_ _04337_ enc_block.round_key\[66\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_87_347 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_213_692 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15664_ VGND VPWR VPWR VGND _10953_ _10508_ _10463_ _11121_ sky130_fd_sc_hd__or3_2
XFILLER_0_198_894 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12876_ VGND VPWR VGND VPWR _07877_ keymem.key_mem\[10\]\[71\] _08405_ _08407_ _08408_
+ _08020_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_73_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_201_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17403_ VPWR VGND VGND VPWR _10327_ _03487_ key[100] sky130_fd_sc_hd__nor2_2
X_14615_ VGND VPWR VGND VPWR _09517_ keymem.prev_key0_reg\[4\] _10080_ _10081_ _10083_
+ sky130_fd_sc_hd__a31o_2
X_11827_ VGND VPWR result[80] _07477_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_5_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18383_ VGND VPWR _04276_ _03977_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15595_ VGND VPWR VGND VPWR _11051_ _11050_ _11053_ _11052_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_28_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17334_ VGND VPWR _03427_ _03426_ VPWR VGND sky130_fd_sc_hd__buf_1
X_11758_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[14\] dec_new_block\[46\]
+ _07443_ sky130_fd_sc_hd__mux2_2
X_14546_ VPWR VGND VGND VPWR _09222_ _10014_ _09029_ sky130_fd_sc_hd__nor2_2
XFILLER_0_172_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17265_ VGND VPWR VPWR VGND _03296_ keymem.key_mem\[14\]\[84\] _03364_ _03365_ sky130_fd_sc_hd__mux2_2
X_14477_ _09086_ _09946_ _09047_ _09945_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_11689_ VGND VPWR result[11] _07408_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_10_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19004_ VGND VPWR VGND VPWR _03959_ block[58] _04834_ _04833_ sky130_fd_sc_hd__a21oi_2
X_16216_ VGND VPWR _02380_ _11236_ _02381_ _11482_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_113_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_148_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13428_ VPWR VGND VPWR VGND _08904_ keymem.key_mem\[12\]\[126\] _07807_ keymem.key_mem\[2\]\[126\]
+ _07698_ _08905_ sky130_fd_sc_hd__a221o_2
X_17196_ VGND VPWR VGND VPWR _03303_ _03302_ _02927_ key[77] sky130_fd_sc_hd__o21a_2
XFILLER_0_84_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16147_ VGND VPWR VGND VPWR _11365_ _11427_ _11344_ _11316_ _11601_ sky130_fd_sc_hd__a2bb2o_2
X_13359_ VGND VPWR VGND VPWR _07835_ keymem.key_mem\[13\]\[119\] _08840_ _08842_ _08843_
+ _08736_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_45_1246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_166_1_Left_433 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_347 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_220_1004 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_126_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16078_ VGND VPWR VGND VPWR _11532_ _11502_ _11533_ _09240_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_121_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_134_2_Left_605 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15029_ VGND VPWR VGND VPWR _10471_ _10479_ _10486_ _10493_ _10492_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_227_228 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19906_ VGND VPWR VPWR VGND _05361_ keymem.key_mem\[11\]\[109\] _03550_ _05365_ sky130_fd_sc_hd__mux2_2
XFILLER_0_196_1537 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19837_ VGND VPWR VPWR VGND _05328_ keymem.key_mem\[11\]\[76\] _03295_ _05329_ sky130_fd_sc_hd__mux2_2
XFILLER_0_209_987 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_732 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19768_ VGND VPWR VPWR VGND _05292_ keymem.key_mem\[11\]\[43\] _02985_ _05293_ sky130_fd_sc_hd__mux2_2
XFILLER_0_155_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_74 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18719_ VGND VPWR _04577_ enc_block.block_w0_reg\[6\] _04372_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_91_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_78_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19699_ VGND VPWR _00638_ _05256_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_155_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21730_ VGND VPWR VPWR VGND _06330_ _03216_ keymem.key_mem\[4\]\[67\] _06335_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_306 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_231_1166 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21661_ VGND VPWR VPWR VGND _06297_ _02893_ keymem.key_mem\[4\]\[34\] _06299_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23400_ VPWR VGND _07272_ _07271_ enc_block.round_key\[19\] VPWR VGND sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_135_2_Right_207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20612_ VGND VPWR VPWR VGND _05736_ _03108_ keymem.key_mem\[8\]\[56\] _05740_ sky130_fd_sc_hd__mux2_2
X_24380_ VGND VPWR VPWR VGND clk _00873_ reset_n keymem.key_mem\[10\]\[117\] sky130_fd_sc_hd__dfrtp_2
X_21592_ VGND VPWR _06262_ _06258_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_778 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_46_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23331_ VPWR VGND VGND VPWR _07192_ _07210_ _04116_ sky130_fd_sc_hd__nor2_2
XFILLER_0_6_330 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20543_ VGND VPWR VPWR VGND _05703_ _02660_ keymem.key_mem\[8\]\[23\] _05704_ sky130_fd_sc_hd__mux2_2
XFILLER_0_7_886 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_104_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_116_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_127_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23262_ VPWR VGND VPWR VGND _07147_ _04874_ _07146_ enc_block.block_w3_reg\[5\] _07115_
+ _02310_ sky130_fd_sc_hd__a221o_2
XFILLER_0_166_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20474_ VGND VPWR _01003_ _05666_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_42_450 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_131_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_601 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_67_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_104_338 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25001_ VGND VPWR VPWR VGND clk _01494_ reset_n keymem.key_mem\[5\]\[98\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_1_Left_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_127_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22213_ VGND VPWR VPWR VGND _06589_ _02903_ keymem.key_mem\[2\]\[35\] _06594_ sky130_fd_sc_hd__mux2_2
XFILLER_0_162_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23193_ VGND VPWR VGND VPWR _02304_ _07084_ _06888_ keymem.prev_key1_reg\[127\] sky130_fd_sc_hd__o21a_2
XFILLER_0_30_634 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_66_2_Left_537 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22144_ VGND VPWR _01782_ _06557_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_238_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1150 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22075_ VGND VPWR VPWR VGND _06516_ _05031_ keymem.key_mem\[3\]\[99\] _06520_ sky130_fd_sc_hd__mux2_2
X_21026_ VGND VPWR _01260_ _05961_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_103_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_946 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25834_ VGND VPWR VPWR VGND clk _02327_ reset_n enc_block.block_w3_reg\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_138_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1356 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25765_ keymem.prev_key1_reg\[81\] clk _02258_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22977_ VGND VPWR VGND VPWR _02219_ _06953_ _06916_ keymem.prev_key1_reg\[42\] sky130_fd_sc_hd__o21a_2
XFILLER_0_173_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_180_2_Left_651 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_74_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12730_ VGND VPWR VGND VPWR _08277_ _07731_ keymem.key_mem\[13\]\[56\] _08274_ _08276_
+ sky130_fd_sc_hd__a211o_2
X_24716_ VGND VPWR VPWR VGND clk _01209_ reset_n keymem.key_mem\[7\]\[69\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21928_ VPWR VGND keymem.key_mem\[3\]\[30\] _06442_ _06439_ VPWR VGND sky130_fd_sc_hd__and2_2
X_25696_ keymem.prev_key1_reg\[12\] clk _02189_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_139_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_38_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_70_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_214_1364 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12661_ VPWR VGND VPWR VGND _08213_ keymem.key_mem\[9\]\[50\] _07717_ keymem.key_mem\[10\]\[50\]
+ _07865_ _08214_ sky130_fd_sc_hd__a221o_2
X_21859_ VGND VPWR _06403_ _06402_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24647_ VGND VPWR VPWR VGND clk _01140_ reset_n keymem.key_mem\[7\]\[0\] sky130_fd_sc_hd__dfrtp_2
X_14400_ VPWR VGND VGND VPWR _09869_ key[131] _09868_ sky130_fd_sc_hd__nand2_2
X_15380_ VGND VPWR _10840_ _10482_ _10841_ _10588_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_12592_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[43\] _07667_ keymem.key_mem\[8\]\[43\]
+ _07540_ _08152_ sky130_fd_sc_hd__a22o_2
X_24578_ VGND VPWR VPWR VGND clk _01071_ reset_n keymem.key_mem\[8\]\[59\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_249_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_1202 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14331_ VGND VPWR VGND VPWR _09204_ _09684_ _09801_ _09125_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_110_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23529_ VGND VPWR VPWR VGND clk _00030_ reset_n keymem.key_mem\[14\]\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_107_143 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14262_ VGND VPWR _09732_ _08927_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17050_ VGND VPWR VGND VPWR _03172_ _03152_ key[190] _03167_ _03171_ sky130_fd_sc_hd__a211o_2
XFILLER_0_145_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_271 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_149_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16001_ VGND VPWR _11456_ _09927_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13213_ VGND VPWR VGND VPWR _07580_ keymem.key_mem\[12\]\[104\] _08707_ _08709_ _08712_
+ _08711_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_46_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_145_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14193_ VPWR VGND VGND VPWR _09125_ _09664_ _09134_ sky130_fd_sc_hd__nor2_2
XFILLER_0_81_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_46_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13144_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[97\] _08577_ _08649_ _08645_ _08650_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_260_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_57_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17952_ VGND VPWR _00248_ _03899_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13075_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[91\] _07779_ keymem.key_mem\[12\]\[91\]
+ _07807_ _08587_ sky130_fd_sc_hd__a22o_2
XFILLER_0_178_1223 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16903_ VGND VPWR VGND VPWR _03038_ _02928_ _02927_ key[49] sky130_fd_sc_hd__o21a_2
XFILLER_0_256_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12026_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[1\] _07535_ _07627_ _07617_ _07628_
+ sky130_fd_sc_hd__o22a_2
X_17883_ VPWR VGND VPWR VGND _03852_ keymem.prev_key1_reg\[86\] sky130_fd_sc_hd__inv_2
XFILLER_0_224_209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_228_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_218_784 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_121_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19622_ VGND VPWR VPWR VGND _05205_ _05041_ keymem.key_mem\[12\]\[104\] _05214_ sky130_fd_sc_hd__mux2_2
X_16834_ _10895_ _02975_ _10894_ _10896_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_73_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19553_ VPWR VGND keymem.key_mem\[12\]\[71\] _05178_ _05173_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_233_776 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_92_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16765_ VPWR VGND VPWR VGND _02912_ _10902_ _02907_ key[164] _02875_ _02913_ sky130_fd_sc_hd__a221o_2
XFILLER_0_152_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13977_ VPWR VGND VPWR VGND _09261_ _09246_ _09315_ _09297_ _09449_ sky130_fd_sc_hd__or4_2
X_18504_ VGND VPWR _04385_ enc_block.block_w0_reg\[6\] _04384_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15716_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[19\] _08954_ _11172_ _08941_ _11170_
+ _11171_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_92_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12928_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[76\] _07632_ keymem.key_mem\[11\]\[76\]
+ _07861_ _08455_ sky130_fd_sc_hd__a22o_2
X_19484_ VGND VPWR _00538_ _05141_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_1083 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_53_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16696_ VGND VPWR _02849_ keymem.prev_key0_reg\[31\] _02848_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_232_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18435_ VGND VPWR _04322_ _04319_ _04321_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15647_ VPWR VGND VGND VPWR _11104_ _10336_ _10359_ sky130_fd_sc_hd__nand2_2
XFILLER_0_28_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12859_ VPWR VGND VPWR VGND _08392_ keymem.key_mem\[3\]\[69\] _08009_ keymem.key_mem\[8\]\[69\]
+ _08265_ _08393_ sky130_fd_sc_hd__a221o_2
XFILLER_0_232_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_222 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_132_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18366_ VPWR VGND VGND VPWR _04261_ _04010_ _04260_ sky130_fd_sc_hd__nand2_2
X_15578_ VGND VPWR VGND VPWR _11037_ _11036_ _11035_ _09866_ _11034_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_22_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17317_ VGND VPWR VGND VPWR _02736_ _02735_ _02708_ _03411_ sky130_fd_sc_hd__a21o_2
XFILLER_0_28_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14529_ VGND VPWR _09643_ _09107_ _09997_ _09174_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_18297_ VPWR VGND VPWR VGND _04198_ block[116] _04076_ enc_block.block_w1_reg\[20\]
+ _04171_ _04199_ sky130_fd_sc_hd__a221o_2
XFILLER_0_22_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17248_ VGND VPWR VPWR VGND _09717_ _02396_ keymem.prev_key0_reg\[83\] _03349_ sky130_fd_sc_hd__or3_2
XFILLER_0_163_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_472 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17179_ VPWR VGND VGND VPWR _03288_ keymem.key_mem\[14\]\[75\] _09541_ sky130_fd_sc_hd__nand2_2
XFILLER_0_51_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20190_ VGND VPWR VPWR VGND _05515_ _03580_ keymem.key_mem\[10\]\[114\] _05516_ sky130_fd_sc_hd__mux2_2
XFILLER_0_121_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_259_1055 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_209_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_710 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_264_890 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_37_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22900_ VGND VPWR VPWR VGND _06878_ _06905_ keymem.prev_key1_reg\[13\] _06906_ sky130_fd_sc_hd__mux2_2
XFILLER_0_236_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23880_ VGND VPWR VPWR VGND clk _00373_ reset_n keymem.key_mem\[13\]\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22831_ VPWR VGND VGND VPWR _06863_ keymem.key_mem_we _06861_ sky130_fd_sc_hd__nand2_2
XFILLER_0_170_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_223_275 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_211_415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_196_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22762_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[77\] _06837_ _06836_ _04995_ _02113_
+ sky130_fd_sc_hd__a22o_2
X_25550_ VGND VPWR VPWR VGND clk _02043_ reset_n keymem.key_mem\[0\]\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_250_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21713_ VGND VPWR VPWR VGND _06319_ _03139_ keymem.key_mem\[4\]\[59\] _06326_ sky130_fd_sc_hd__mux2_2
X_24501_ VGND VPWR VPWR VGND clk _00994_ reset_n keymem.key_mem\[9\]\[110\] sky130_fd_sc_hd__dfrtp_2
X_25481_ VGND VPWR VPWR VGND clk _01974_ reset_n keymem.key_mem\[1\]\[66\] sky130_fd_sc_hd__dfrtp_2
X_22693_ VGND VPWR _02071_ _06817_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_13_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24432_ VGND VPWR VPWR VGND clk _00925_ reset_n keymem.key_mem\[9\]\[41\] sky130_fd_sc_hd__dfrtp_2
X_21644_ VGND VPWR VPWR VGND _06286_ _02742_ keymem.key_mem\[4\]\[26\] _06290_ sky130_fd_sc_hd__mux2_2
XFILLER_0_19_255 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_136_2_Right_208 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24363_ VGND VPWR VPWR VGND clk _00856_ reset_n keymem.key_mem\[10\]\[100\] sky130_fd_sc_hd__dfrtp_2
X_21575_ VGND VPWR VPWR VGND _06242_ _03640_ keymem.key_mem\[5\]\[123\] _06252_ sky130_fd_sc_hd__mux2_2
XFILLER_0_19_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_394 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23314_ VPWR VGND _07194_ _07128_ enc_block.block_w2_reg\[2\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_209_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20526_ VGND VPWR VPWR VGND _05692_ _11148_ keymem.key_mem\[8\]\[15\] _05695_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24294_ VGND VPWR VPWR VGND clk _00787_ reset_n keymem.key_mem\[10\]\[31\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_144_271 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_182 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_166_1171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_43_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23245_ VGND VPWR _07132_ _07130_ _07131_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_1110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20457_ VGND VPWR _00995_ _05657_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_28_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23176_ VGND VPWR VGND VPWR _03623_ _03622_ _03626_ _07074_ sky130_fd_sc_hd__a21o_2
XFILLER_0_28_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20388_ VGND VPWR _00962_ _05621_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_63_1187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_526 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22127_ VGND VPWR VPWR VGND _06538_ _05083_ keymem.key_mem\[3\]\[124\] _06547_ sky130_fd_sc_hd__mux2_2
XFILLER_0_24_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22058_ VPWR VGND keymem.key_mem\[3\]\[91\] _06511_ _06405_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_265_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13900_ VPWR VGND VGND VPWR _09372_ _09370_ _09371_ sky130_fd_sc_hd__nand2_2
X_21009_ VGND VPWR _01252_ _05952_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14880_ VPWR VGND VPWR VGND _10339_ _10344_ _10345_ _09192_ _10337_ sky130_fd_sc_hd__or4b_2
XFILLER_0_216_1415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13831_ VGND VPWR _09303_ _09297_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25817_ VGND VPWR VPWR VGND clk _02310_ reset_n enc_block.block_w3_reg\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_214_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_138_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_189_1_Right_790 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16550_ VGND VPWR VGND VPWR _02694_ _02693_ keymem.prev_key1_reg\[121\] _02709_ sky130_fd_sc_hd__a21o_2
XFILLER_0_138_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13762_ VPWR VGND VGND VPWR _09134_ _09234_ _09148_ sky130_fd_sc_hd__nor2_2
X_25748_ keymem.prev_key1_reg\[64\] clk _02241_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_230_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_74_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15501_ VPWR VGND _10948_ _10961_ _10960_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_211_960 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12713_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[55\] _07918_ keymem.key_mem\[12\]\[55\]
+ _07806_ _08261_ sky130_fd_sc_hd__a22o_2
X_16481_ VGND VPWR _02642_ keymem.prev_key0_reg\[55\] keymem.prev_key0_reg\[87\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
X_13693_ VGND VPWR VGND VPWR _09075_ _09093_ _09119_ _09165_ _09164_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_69_199 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_214_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_210_1014 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25679_ VGND VPWR VPWR VGND clk _02172_ reset_n keymem.round_ctr_reg\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18220_ VPWR VGND _04128_ enc_block.block_w3_reg\[6\] enc_block.block_w3_reg\[5\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_15432_ _10861_ _10893_ keymem.round_ctr_reg\[0\] _10892_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_210_492 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12644_ VPWR VGND VPWR VGND _08198_ keymem.key_mem\[6\]\[48\] _07711_ keymem.key_mem\[1\]\[48\]
+ _07671_ _08199_ sky130_fd_sc_hd__a221o_2
XFILLER_0_72_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_127_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18151_ VGND VPWR _04065_ _04064_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12575_ VGND VPWR VGND VPWR _08136_ _07648_ keymem.key_mem\[2\]\[42\] _08135_ _07896_
+ sky130_fd_sc_hd__a211o_2
X_15363_ VGND VPWR _10824_ keymem.prev_key0_reg\[10\] _10825_ _10822_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_25_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17102_ VGND VPWR _00079_ _03218_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_230_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14314_ VPWR VGND VPWR VGND _09784_ _09559_ _09301_ sky130_fd_sc_hd__or2_2
X_18082_ VPWR VGND VPWR VGND _04001_ block[98] _03980_ enc_block.block_w3_reg\[2\]
+ _03978_ _04002_ sky130_fd_sc_hd__a221o_2
XFILLER_0_13_409 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15294_ VPWR VGND VPWR VGND _10756_ _10619_ _10672_ _10572_ _10750_ _10755_ sky130_fd_sc_hd__o311a_2
XFILLER_0_145_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17033_ VPWR VGND VPWR VGND _03156_ keymem.prev_key1_reg\[61\] sky130_fd_sc_hd__inv_2
X_14245_ VGND VPWR VGND VPWR _09714_ _09713_ _09716_ _09715_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_145_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14176_ VGND VPWR VGND VPWR _09067_ _09646_ _09204_ _09050_ _09647_ sky130_fd_sc_hd__o22a_2
XFILLER_0_106_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_46_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13127_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[96\] _07667_ keymem.key_mem\[2\]\[96\]
+ _07732_ _08634_ sky130_fd_sc_hd__a22o_2
X_18984_ VPWR VGND VGND VPWR _04816_ _04591_ _04815_ sky130_fd_sc_hd__nand2_2
XFILLER_0_265_654 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_221_1165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17935_ VGND VPWR VPWR VGND _03874_ _03887_ keymem.prev_key0_reg\[102\] _03888_ sky130_fd_sc_hd__mux2_2
X_13058_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[89\] _08216_ keymem.key_mem\[12\]\[89\]
+ _07722_ _08572_ sky130_fd_sc_hd__a22o_2
XFILLER_0_84_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_721 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12009_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[1\] _07561_ keymem.key_mem\[4\]\[1\]
+ _07551_ _07611_ sky130_fd_sc_hd__a22o_2
XFILLER_0_264_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17866_ VGND VPWR VPWR VGND _03836_ _03840_ keymem.prev_key0_reg\[80\] _03841_ sky130_fd_sc_hd__mux2_2
XFILLER_0_191_1220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19605_ VGND VPWR _05205_ _05091_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_221_702 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16817_ VPWR VGND VPWR VGND _02960_ _02864_ _10664_ _02957_ _02959_ _02866_ sky130_fd_sc_hd__o311a_2
XFILLER_0_156_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17797_ VGND VPWR _03794_ _09638_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_255_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_735 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19536_ VPWR VGND keymem.key_mem\[12\]\[63\] _05169_ _05158_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_156_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16748_ VPWR VGND VPWR VGND _02897_ keymem.prev_key1_reg\[35\] sky130_fd_sc_hd__inv_2
XFILLER_0_117_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19467_ VPWR VGND keymem.key_mem\[12\]\[31\] _05132_ _05128_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_5_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16679_ VPWR VGND _02833_ keymem.prev_key1_reg\[62\] keymem.prev_key1_reg\[30\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_14_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18418_ VPWR VGND _04306_ enc_block.block_w2_reg\[16\] enc_block.block_w3_reg\[8\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_57_862 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_63_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_88_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19398_ VPWR VGND VPWR VGND _05094_ _09538_ _08925_ sky130_fd_sc_hd__or2_2
X_18349_ VPWR VGND VPWR VGND _04245_ block[121] _04213_ enc_block.block_w0_reg\[25\]
+ _04171_ _04246_ sky130_fd_sc_hd__a221o_2
XFILLER_0_267_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_394 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21360_ VGND VPWR _01416_ _06139_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_1105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_163_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20311_ VGND VPWR _00925_ _05581_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_167_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21291_ VGND VPWR VPWR VGND _06098_ _03600_ keymem.key_mem\[6\]\[117\] _06102_ sky130_fd_sc_hd__mux2_2
XFILLER_0_128_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_263 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23030_ VGND VPWR _02241_ _06984_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20242_ VGND VPWR VPWR VGND _05535_ _10747_ keymem.key_mem\[9\]\[9\] _05545_ sky130_fd_sc_hd__mux2_2
XFILLER_0_124_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_857 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20173_ VGND VPWR VPWR VGND _05504_ _03533_ keymem.key_mem\[10\]\[106\] _05507_ sky130_fd_sc_hd__mux2_2
XFILLER_0_25_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24981_ VGND VPWR VPWR VGND clk _01474_ reset_n keymem.key_mem\[5\]\[78\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_1142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_239_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23932_ VGND VPWR VPWR VGND clk _00425_ reset_n keymem.key_mem\[13\]\[53\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_174_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23863_ VGND VPWR VPWR VGND clk _00356_ reset_n enc_block.block_w2_reg\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_139_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25602_ VGND VPWR VPWR VGND clk _02095_ reset_n keymem.key_mem\[0\]\[59\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_36_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22814_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[113\] _06860_ _06859_ _05060_ _02149_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_170_1326 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23794_ VGND VPWR VPWR VGND clk _00287_ reset_n enc_block.block_w0_reg\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_71_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25533_ VGND VPWR VPWR VGND clk _02026_ reset_n keymem.key_mem\[1\]\[118\] sky130_fd_sc_hd__dfrtp_2
X_22745_ VGND VPWR VPWR VGND _06833_ keymem.key_mem\[0\]\[67\] _03217_ _06838_ sky130_fd_sc_hd__mux2_2
XFILLER_0_215_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_211_1345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_181_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_133_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25464_ VGND VPWR VPWR VGND clk _01957_ reset_n keymem.key_mem\[1\]\[49\] sky130_fd_sc_hd__dfrtp_2
X_22676_ VGND VPWR VPWR VGND _06809_ keymem.key_mem\[0\]\[26\] _02743_ _06810_ sky130_fd_sc_hd__mux2_2
XFILLER_0_211_1356 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_512 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_63_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_1142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24415_ VGND VPWR VPWR VGND clk _00908_ reset_n keymem.key_mem\[9\]\[24\] sky130_fd_sc_hd__dfrtp_2
X_21627_ VGND VPWR VPWR VGND _06275_ _02339_ keymem.key_mem\[4\]\[18\] _06281_ sky130_fd_sc_hd__mux2_2
X_25395_ VGND VPWR VPWR VGND clk _01888_ reset_n keymem.key_mem\[2\]\[108\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_8_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_556 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_137_2_Right_209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_707 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12360_ VPWR VGND VPWR VGND _07940_ keymem.key_mem\[4\]\[22\] _07637_ keymem.key_mem\[2\]\[22\]
+ _07546_ _07941_ sky130_fd_sc_hd__a221o_2
XFILLER_0_168_1277 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24346_ VGND VPWR VPWR VGND clk _00839_ reset_n keymem.key_mem\[10\]\[83\] sky130_fd_sc_hd__dfrtp_2
X_21558_ VGND VPWR _01510_ _06243_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_23_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20509_ VGND VPWR VPWR VGND _05680_ _10369_ keymem.key_mem\[8\]\[7\] _05686_ sky130_fd_sc_hd__mux2_2
X_12291_ VGND VPWR _07877_ _07876_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24277_ VGND VPWR VPWR VGND clk _00770_ reset_n keymem.key_mem\[10\]\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_107_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21489_ VGND VPWR VPWR VGND _06196_ _03346_ keymem.key_mem\[5\]\[82\] _06207_ sky130_fd_sc_hd__mux2_2
XFILLER_0_146_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14030_ VGND VPWR VPWR VGND _09343_ _09366_ _09362_ _09502_ sky130_fd_sc_hd__or3_2
X_23228_ VGND VPWR _07116_ enc_block.block_w3_reg\[31\] enc_block.block_w1_reg\[11\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_82_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1093 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23159_ VGND VPWR VGND VPWR _07064_ _03575_ _06890_ _06924_ _03579_ sky130_fd_sc_hd__a211o_2
XFILLER_0_38_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15981_ VPWR VGND VPWR VGND _11424_ _11436_ _11431_ _11415_ _11437_ sky130_fd_sc_hd__or4_2
XFILLER_0_59_1009 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_257_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17720_ VPWR VGND VPWR VGND _02784_ _03746_ keymem.prev_key0_reg\[28\] _03730_ _00169_
+ sky130_fd_sc_hd__a22o_2
X_14932_ VPWR VGND VPWR VGND _10396_ enc_block.block_w0_reg\[8\] _09273_ sky130_fd_sc_hd__or2_2
XFILLER_0_262_657 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17651_ VGND VPWR VPWR VGND _03681_ _03696_ keymem.prev_key0_reg\[9\] _03697_ sky130_fd_sc_hd__mux2_2
X_14863_ VGND VPWR _10328_ _09512_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_243_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_199_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16602_ VGND VPWR _02759_ keymem.prev_key1_reg\[27\] keymem.prev_key1_reg\[59\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
X_13814_ VGND VPWR VGND VPWR _09286_ enc_block.block_w2_reg\[28\] enc_block.sword_ctr_reg\[1\]
+ enc_block.sword_ctr_reg\[0\] sky130_fd_sc_hd__and3b_2
XFILLER_0_153_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1256 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17582_ VPWR VGND VGND VPWR _03642_ _03240_ _02771_ sky130_fd_sc_hd__nand2_2
X_14794_ VGND VPWR VGND VPWR _09917_ _10260_ _10255_ _10259_ _10250_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_114_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19321_ VPWR VGND keymem.key_mem_we _05041_ _03518_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_97_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16533_ VPWR VGND VPWR VGND _02692_ keymem.rcon_logic.tmp_rcon\[2\] sky130_fd_sc_hd__inv_2
X_13745_ VPWR VGND VPWR VGND _08963_ _09027_ _09017_ _08957_ _09217_ sky130_fd_sc_hd__or4_2
XFILLER_0_225_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_175_1_Left_442 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19252_ VGND VPWR VPWR VGND _04993_ _04997_ keymem.key_mem\[13\]\[78\] _04998_ sky130_fd_sc_hd__mux2_2
X_16464_ VGND VPWR VGND VPWR _02624_ _02623_ _02625_ _02622_ _02621_ sky130_fd_sc_hd__nand4_2
X_13676_ VGND VPWR _09148_ _09147_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_155_322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_143_2_Left_614 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18203_ VPWR VGND VGND VPWR _04112_ _04113_ _04077_ sky130_fd_sc_hd__nor2_2
X_15415_ VGND VPWR VGND VPWR _10751_ _10489_ _10876_ _10595_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_241_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_72_128 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12627_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[47\] _07845_ keymem.key_mem\[12\]\[47\]
+ _07788_ _08183_ sky130_fd_sc_hd__a22o_2
X_19183_ VGND VPWR _00422_ _04956_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_182_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16395_ _11461_ _02557_ _11285_ _11462_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_26_545 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18134_ VPWR VGND VPWR VGND _04049_ block[102] _03980_ enc_block.block_w3_reg\[6\]
+ _04007_ _04050_ sky130_fd_sc_hd__a221o_2
X_15346_ VPWR VGND VGND VPWR _10414_ _10458_ _10808_ _10557_ _10469_ sky130_fd_sc_hd__o22ai_2
X_12558_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[40\] _07748_ keymem.key_mem\[9\]\[40\]
+ _07705_ _08121_ sky130_fd_sc_hd__a22o_2
XFILLER_0_26_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18065_ VGND VPWR _03986_ _03984_ _03985_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_227_1374 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15277_ VGND VPWR VPWR VGND _10740_ keymem.prev_key1_reg\[73\] _10737_ _10738_ _08927_
+ sky130_fd_sc_hd__o31a_2
X_12489_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[34\] _07659_ keymem.key_mem\[1\]\[34\]
+ _07714_ _08058_ sky130_fd_sc_hd__a22o_2
XFILLER_0_1_623 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17016_ VGND VPWR VPWR VGND _03084_ keymem.key_mem\[14\]\[59\] _03140_ _03141_ sky130_fd_sc_hd__mux2_2
X_14228_ VGND VPWR VGND VPWR _09698_ _09057_ _09087_ _09062_ _09699_ sky130_fd_sc_hd__a31o_2
XFILLER_0_240_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14159_ VGND VPWR VGND VPWR _09629_ _09589_ keymem.prev_key1_reg\[97\] _09630_ sky130_fd_sc_hd__a21o_2
XFILLER_0_10_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18967_ VGND VPWR _04801_ enc_block.block_w3_reg\[21\] enc_block.block_w2_reg\[30\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_201_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17918_ VGND VPWR _03876_ _03211_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18898_ VPWR VGND VGND VPWR _04739_ _04736_ _04737_ sky130_fd_sc_hd__nand2_2
X_17849_ VGND VPWR VPWR VGND _03812_ key[203] keymem.prev_key1_reg\[75\] _03829_ sky130_fd_sc_hd__mux2_2
X_20860_ VGND VPWR VPWR VGND _05867_ _04939_ keymem.key_mem\[7\]\[42\] _05874_ sky130_fd_sc_hd__mux2_2
XFILLER_0_221_565 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_53_1131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19519_ VGND VPWR VPWR VGND _05151_ _04963_ keymem.key_mem\[12\]\[55\] _05160_ sky130_fd_sc_hd__mux2_2
X_20791_ VGND VPWR VGND VPWR _05836_ keymem.key_mem_we _10836_ _05821_ _01150_ sky130_fd_sc_hd__a31o_2
XFILLER_0_18_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_2_Left_546 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_48_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_202_790 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_723 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22530_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[65\] _06737_ _06736_ _04975_ _01973_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_48_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_64_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_88_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22461_ VGND VPWR _01932_ _06724_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_130_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24200_ VGND VPWR VPWR VGND clk _00693_ reset_n keymem.key_mem\[11\]\[65\] sky130_fd_sc_hd__dfrtp_2
X_21412_ VGND VPWR VPWR VGND _06162_ _03006_ keymem.key_mem\[5\]\[45\] _06167_ sky130_fd_sc_hd__mux2_2
XFILLER_0_161_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_95 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25180_ VGND VPWR VPWR VGND clk _01673_ reset_n keymem.key_mem\[3\]\[21\] sky130_fd_sc_hd__dfrtp_2
X_22392_ VGND VPWR _01900_ _06687_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_32_515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24131_ VGND VPWR VPWR VGND clk _00624_ reset_n keymem.key_mem\[12\]\[124\] sky130_fd_sc_hd__dfrtp_2
X_21343_ VGND VPWR VPWR VGND _06128_ _10976_ keymem.key_mem\[5\]\[12\] _06131_ sky130_fd_sc_hd__mux2_2
XFILLER_0_128_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24062_ VGND VPWR VPWR VGND clk _00555_ reset_n keymem.key_mem\[12\]\[55\] sky130_fd_sc_hd__dfrtp_2
X_21274_ VGND VPWR VPWR VGND _06087_ _03550_ keymem.key_mem\[6\]\[109\] _06093_ sky130_fd_sc_hd__mux2_2
XFILLER_0_25_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23013_ VPWR VGND VPWR VGND _06975_ keymem.prev_key1_reg\[57\] _06926_ sky130_fd_sc_hd__or2_2
X_20225_ VGND VPWR _00884_ _05536_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_99_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_816 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_200_1024 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20156_ VGND VPWR VPWR VGND _05493_ _03480_ keymem.key_mem\[10\]\[98\] _05498_ sky130_fd_sc_hd__mux2_2
XFILLER_0_99_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20087_ VGND VPWR VPWR VGND _05457_ _03202_ keymem.key_mem\[10\]\[65\] _05462_ sky130_fd_sc_hd__mux2_2
X_24964_ VGND VPWR VPWR VGND clk _01457_ reset_n keymem.key_mem\[5\]\[61\] sky130_fd_sc_hd__dfrtp_2
X_23915_ VGND VPWR VPWR VGND clk _00408_ reset_n keymem.key_mem\[13\]\[36\] sky130_fd_sc_hd__dfrtp_2
X_24895_ VGND VPWR VPWR VGND clk _01388_ reset_n keymem.key_mem\[6\]\[120\] sky130_fd_sc_hd__dfrtp_2
X_11860_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[1\] dec_new_block\[97\]
+ _07494_ sky130_fd_sc_hd__mux2_2
X_23846_ VGND VPWR VPWR VGND clk _00339_ reset_n enc_block.block_w1_reg\[31\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_86_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_170_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_778 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11791_ VGND VPWR result[62] _07459_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20989_ VGND VPWR VPWR VGND _05934_ _05039_ keymem.key_mem\[7\]\[103\] _05942_ sky130_fd_sc_hd__mux2_2
XFILLER_0_212_598 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23777_ VGND VPWR VPWR VGND clk _00270_ reset_n enc_block.round\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_36_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13530_ VGND VPWR _09002_ _08941_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25516_ VGND VPWR VPWR VGND clk _02009_ reset_n keymem.key_mem\[1\]\[101\] sky130_fd_sc_hd__dfrtp_2
X_22728_ VGND VPWR VPWR VGND _06822_ keymem.key_mem\[0\]\[59\] _03140_ _06829_ sky130_fd_sc_hd__mux2_2
XFILLER_0_149_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_94_286 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25447_ VGND VPWR VPWR VGND clk _01940_ reset_n keymem.key_mem\[1\]\[32\] sky130_fd_sc_hd__dfrtp_2
X_13461_ VPWR VGND VGND VPWR keymem.round_ctr_reg\[3\] _08933_ keymem.round_ctr_reg\[2\]
+ sky130_fd_sc_hd__nor2_2
XFILLER_0_246_1205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22659_ VGND VPWR VPWR VGND _06798_ keymem.key_mem\[0\]\[18\] _02340_ _06801_ sky130_fd_sc_hd__mux2_2
XFILLER_0_152_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15200_ VGND VPWR _00020_ _10663_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12412_ VGND VPWR VGND VPWR _07984_ keymem.key_mem\[14\]\[27\] _07985_ _07987_ _07988_
+ _07662_ sky130_fd_sc_hd__a2111o_2
X_16180_ VGND VPWR VGND VPWR _11292_ _11389_ _11271_ _02345_ sky130_fd_sc_hd__a21o_2
XFILLER_0_63_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25378_ VGND VPWR VPWR VGND clk _01871_ reset_n keymem.key_mem\[2\]\[91\] sky130_fd_sc_hd__dfrtp_2
X_13392_ VPWR VGND VPWR VGND _08872_ keymem.key_mem\[13\]\[122\] _08125_ keymem.key_mem\[11\]\[122\]
+ _07902_ _08873_ sky130_fd_sc_hd__a221o_2
XFILLER_0_152_358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15131_ VGND VPWR _10595_ _10594_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24329_ VGND VPWR VPWR VGND clk _00822_ reset_n keymem.key_mem\[10\]\[66\] sky130_fd_sc_hd__dfrtp_2
X_12343_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[21\] _07618_ keymem.key_mem\[6\]\[21\]
+ _07759_ _07925_ sky130_fd_sc_hd__a22o_2
XFILLER_0_209_1060 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_107_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15062_ VPWR VGND VPWR VGND _10483_ _10466_ _10453_ _10439_ _10526_ sky130_fd_sc_hd__or4_2
X_12274_ VGND VPWR _07861_ _07599_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_142_1214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14013_ VPWR VGND VPWR VGND _09260_ _09316_ _09266_ _09253_ _09485_ sky130_fd_sc_hd__or4_2
XFILLER_0_107_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19870_ VGND VPWR VPWR VGND _05339_ keymem.key_mem\[11\]\[92\] _03435_ _05346_ sky130_fd_sc_hd__mux2_2
X_18821_ VGND VPWR _04670_ _04667_ _04669_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18752_ VGND VPWR _04607_ _04605_ _04606_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15964_ VGND VPWR _11420_ _11419_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_263_988 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_257_1378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17703_ VGND VPWR VGND VPWR _03732_ keymem.prev_key1_reg\[24\] _03734_ _03733_ sky130_fd_sc_hd__a21oi_2
X_14915_ VGND VPWR VPWR VGND _10379_ keymem.prev_key1_reg\[72\] _10373_ _10374_ _10378_
+ sky130_fd_sc_hd__o31a_2
X_18683_ VPWR VGND VGND VPWR _04545_ _04319_ _04544_ sky130_fd_sc_hd__nand2_2
X_15895_ VPWR VGND VPWR VGND _11272_ _11208_ _11197_ _11187_ _11351_ sky130_fd_sc_hd__or4_2
XFILLER_0_234_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17634_ VGND VPWR VGND VPWR _10093_ keymem.prev_key1_reg\[4\] _03685_ _03670_ sky130_fd_sc_hd__a21bo_2
X_14846_ _10309_ _10311_ _10308_ _10310_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_81_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17565_ VGND VPWR VPWR VGND _03593_ keymem.key_mem\[14\]\[121\] _03627_ _03628_ sky130_fd_sc_hd__mux2_2
XFILLER_0_203_587 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14777_ VPWR VGND VGND VPWR _10233_ _10243_ _10242_ _10235_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_230_384 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_58_445 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11989_ VGND VPWR _07592_ _07591_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19304_ VGND VPWR VPWR VGND _05025_ _05029_ keymem.key_mem\[13\]\[98\] _05030_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_201_Right_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_46_607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16516_ VGND VPWR VPWR VGND _11109_ _02675_ key[24] _02676_ sky130_fd_sc_hd__mux2_2
XFILLER_0_14_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13728_ VPWR VGND VPWR VGND _09058_ _09039_ _09051_ _09009_ _09200_ sky130_fd_sc_hd__or4_2
XFILLER_0_89_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17496_ VGND VPWR VPWR VGND _03534_ keymem.key_mem\[14\]\[112\] _03567_ _03568_ sky130_fd_sc_hd__mux2_2
XFILLER_0_128_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_821 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19235_ VGND VPWR VPWR VGND _04951_ _04986_ keymem.key_mem\[13\]\[72\] _04987_ sky130_fd_sc_hd__mux2_2
XFILLER_0_14_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16447_ VGND VPWR VPWR VGND _11041_ keymem.key_mem\[14\]\[22\] _02608_ _02609_ sky130_fd_sc_hd__mux2_2
X_13659_ VPWR VGND VGND VPWR _09125_ _09100_ _09053_ _09122_ _09131_ _09130_ sky130_fd_sc_hd__o221a_2
XFILLER_0_128_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19166_ VPWR VGND keymem.key_mem_we _04945_ _03006_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16378_ VGND VPWR _02541_ keymem.prev_key0_reg\[53\] keymem.prev_key0_reg\[85\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18117_ VGND VPWR _04034_ enc_block.block_w0_reg\[29\] _04033_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_186_1196 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15329_ VGND VPWR VGND VPWR _10588_ _10563_ _10584_ _10751_ _10791_ sky130_fd_sc_hd__a31o_2
X_19097_ VGND VPWR _04903_ _04879_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_30_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18048_ VGND VPWR _03970_ _08940_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_125_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_760 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20010_ VGND VPWR _00784_ _05421_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_238_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_94 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_96_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19999_ VGND VPWR VPWR VGND _05413_ _02661_ keymem.key_mem\[10\]\[23\] _05416_ sky130_fd_sc_hd__mux2_2
XFILLER_0_20_1141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_236_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1145 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21961_ VGND VPWR _01697_ _06459_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_213_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_146_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23700_ keymem.prev_key0_reg\[56\] clk _00197_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_55_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_94_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20912_ VGND VPWR VPWR VGND _05880_ _04977_ keymem.key_mem\[7\]\[66\] _05902_ sky130_fd_sc_hd__mux2_2
X_24680_ VGND VPWR VPWR VGND clk _01173_ reset_n keymem.key_mem\[7\]\[33\] sky130_fd_sc_hd__dfrtp_2
X_21892_ VGND VPWR VGND VPWR _06422_ keymem.key_mem_we _11040_ _06420_ _01665_ sky130_fd_sc_hd__a31o_2
XFILLER_0_136_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20843_ VPWR VGND keymem.key_mem\[7\]\[34\] _05865_ _05856_ VPWR VGND sky130_fd_sc_hd__and2_2
X_23631_ VGND VPWR VPWR VGND clk _00132_ reset_n keymem.key_mem\[14\]\[120\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1057 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_178_288 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23562_ VGND VPWR VPWR VGND clk _00063_ reset_n keymem.key_mem\[14\]\[51\] sky130_fd_sc_hd__dfrtp_2
X_20774_ VGND VPWR VGND VPWR _05827_ keymem.key_mem_we _09862_ _05821_ _01142_ sky130_fd_sc_hd__a31o_2
XFILLER_0_71_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25301_ VGND VPWR VPWR VGND clk _01794_ reset_n keymem.key_mem\[2\]\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_193_269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22513_ VGND VPWR VPWR VGND _06739_ keymem.key_mem\[1\]\[57\] _03119_ _06744_ sky130_fd_sc_hd__mux2_2
XFILLER_0_146_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_843 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23493_ VGND VPWR VGND VPWR _03959_ block[30] _07354_ _07353_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_247_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_597 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_342 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_91_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_802 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25232_ VGND VPWR VPWR VGND clk _01725_ reset_n keymem.key_mem\[3\]\[73\] sky130_fd_sc_hd__dfrtp_2
X_22444_ VGND VPWR VPWR VGND _06715_ keymem.key_mem\[1\]\[16\] _11447_ _06716_ sky130_fd_sc_hd__mux2_2
XFILLER_0_45_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_208_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22375_ VGND VPWR _01892_ _06678_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25163_ VGND VPWR VPWR VGND clk _01656_ reset_n keymem.key_mem\[3\]\[4\] sky130_fd_sc_hd__dfrtp_2
X_24114_ VGND VPWR VPWR VGND clk _00607_ reset_n keymem.key_mem\[12\]\[107\] sky130_fd_sc_hd__dfrtp_2
X_21326_ VGND VPWR VPWR VGND _06117_ _10098_ keymem.key_mem\[5\]\[4\] _06122_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_280 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25094_ VGND VPWR VPWR VGND clk _01587_ reset_n keymem.key_mem\[4\]\[63\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_182_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_104_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21257_ VGND VPWR VPWR VGND _06076_ _03499_ keymem.key_mem\[6\]\[101\] _06084_ sky130_fd_sc_hd__mux2_2
X_24045_ VGND VPWR VPWR VGND clk _00538_ reset_n keymem.key_mem\[12\]\[38\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_257_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20208_ VGND VPWR VPWR VGND _05515_ _03640_ keymem.key_mem\[10\]\[123\] _05525_ sky130_fd_sc_hd__mux2_2
X_21188_ VPWR VGND VGND VPWR _06048_ keymem.key_mem\[6\]\[68\] _05985_ sky130_fd_sc_hd__nand2_2
XFILLER_0_141_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20139_ VGND VPWR VPWR VGND _05482_ _03418_ keymem.key_mem\[10\]\[90\] _05489_ sky130_fd_sc_hd__mux2_2
XFILLER_0_102_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_245_988 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24947_ VGND VPWR VPWR VGND clk _01440_ reset_n keymem.key_mem\[5\]\[44\] sky130_fd_sc_hd__dfrtp_2
X_12961_ VGND VPWR VGND VPWR _08485_ _07712_ keymem.key_mem\[6\]\[79\] _08482_ _08484_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_239_1097 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_176_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14700_ VPWR VGND VGND VPWR _09070_ _10167_ _09176_ sky130_fd_sc_hd__nor2_2
XFILLER_0_213_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11912_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[27\] dec_new_block\[123\]
+ _07520_ sky130_fd_sc_hd__mux2_2
X_15680_ VGND VPWR VGND VPWR _10583_ _10536_ _10572_ _10867_ _11137_ sky130_fd_sc_hd__a31o_2
X_12892_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[73\] _07725_ keymem.key_mem\[4\]\[73\]
+ _07854_ _08422_ sky130_fd_sc_hd__a22o_2
X_24878_ VGND VPWR VPWR VGND clk _01371_ reset_n keymem.key_mem\[6\]\[103\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_73_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14631_ VGND VPWR _10099_ _10098_ VPWR VGND sky130_fd_sc_hd__buf_1
X_11843_ VGND VPWR result[88] _07485_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23829_ VGND VPWR VPWR VGND clk _00322_ reset_n enc_block.block_w1_reg\[14\] sky130_fd_sc_hd__dfrtp_2
X_17350_ VPWR VGND VPWR VGND _03441_ key[93] _11543_ sky130_fd_sc_hd__or2_2
X_14562_ VPWR VGND VPWR VGND _09812_ _10029_ _09802_ _09699_ _10030_ sky130_fd_sc_hd__or4_2
X_11774_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[22\] dec_new_block\[54\]
+ _07451_ sky130_fd_sc_hd__mux2_2
XFILLER_0_55_415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16301_ _02463_ _02465_ keymem.prev_key0_reg\[20\] _02464_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_13513_ VGND VPWR _08985_ _08947_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_55_437 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17281_ VGND VPWR VGND VPWR _03379_ _03302_ _02927_ key[86] sky130_fd_sc_hd__o21a_2
X_14493_ VGND VPWR VGND VPWR _09154_ _09095_ _09962_ _09211_ sky130_fd_sc_hd__a21oi_2
X_19020_ VPWR VGND VGND VPWR _04848_ _04637_ _04847_ sky130_fd_sc_hd__nand2_2
X_16232_ VPWR VGND VGND VPWR _02397_ _10189_ _02396_ sky130_fd_sc_hd__nand2_2
X_13444_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[127\] _08027_ _08919_ _08915_ _08920_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_42_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_64_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16163_ VPWR VGND VPWR VGND _11610_ _11616_ _11615_ _11374_ _11617_ sky130_fd_sc_hd__or4_2
XFILLER_0_152_166 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13375_ VGND VPWR enc_block.round_key\[120\] _08857_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15114_ VPWR VGND VGND VPWR _10568_ _10578_ _10496_ sky130_fd_sc_hd__nor2_2
XFILLER_0_50_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12326_ VGND VPWR _07909_ _07742_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_80_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16094_ VGND VPWR _00029_ _11548_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_84_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15045_ VPWR VGND VPWR VGND _10483_ _10409_ _10403_ _10412_ _10509_ sky130_fd_sc_hd__or4_2
XFILLER_0_50_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19922_ VGND VPWR _00744_ _05373_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_2_Left_270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12257_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[14\] _07845_ keymem.key_mem\[3\]\[14\]
+ _07844_ _07846_ sky130_fd_sc_hd__a22o_2
XFILLER_0_76_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1152 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_236_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19853_ VGND VPWR VPWR VGND _05328_ keymem.key_mem\[11\]\[84\] _03364_ _05337_ sky130_fd_sc_hd__mux2_2
X_12188_ VGND VPWR _07781_ _07658_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_120_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18804_ VPWR VGND VGND VPWR _04654_ _04655_ _04042_ sky130_fd_sc_hd__nor2_2
XFILLER_0_120_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19784_ VGND VPWR VPWR VGND _05292_ keymem.key_mem\[11\]\[51\] _03068_ _05301_ sky130_fd_sc_hd__mux2_2
X_16996_ VPWR VGND VPWR VGND _03122_ key[58] _09719_ sky130_fd_sc_hd__or2_2
XFILLER_0_247_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18735_ VGND VPWR _04591_ enc_block.block_w2_reg\[31\] enc_block.block_w0_reg\[8\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15947_ VPWR VGND VPWR VGND _11227_ _11273_ _11289_ _11225_ _11403_ sky130_fd_sc_hd__or4_2
XFILLER_0_251_947 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_194_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_162_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18666_ VPWR VGND VPWR VGND _04530_ _04461_ _04529_ sky130_fd_sc_hd__or2_2
X_15878_ VPWR VGND VPWR VGND _11173_ _11248_ _11180_ _11166_ _11334_ sky130_fd_sc_hd__or4_2
XFILLER_0_91_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14829_ VPWR VGND VGND VPWR _10293_ _10294_ _09368_ sky130_fd_sc_hd__nor2_2
X_17617_ VPWR VGND VGND VPWR _03672_ keymem.key_mem_we reset_n sky130_fd_sc_hd__nand2_2
X_18597_ VGND VPWR _04468_ _04159_ _00324_ _04317_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_263_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17548_ VPWR VGND VPWR VGND _03612_ _03494_ _03609_ key[247] _03527_ _03613_ sky130_fd_sc_hd__a221o_2
XFILLER_0_89_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_128_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_131_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17479_ VPWR VGND VPWR VGND _03553_ key[110] _09987_ sky130_fd_sc_hd__or2_2
XFILLER_0_41_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19218_ VGND VPWR _00437_ _04976_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_27_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20490_ VGND VPWR _01011_ _05674_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_143_122 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_138_1_Left_405 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_846 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19149_ VGND VPWR VPWR VGND _04928_ _04933_ keymem.key_mem\[13\]\[39\] _04934_ sky130_fd_sc_hd__mux2_2
XFILLER_0_15_868 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22160_ VGND VPWR VPWR VGND _06565_ _10835_ keymem.key_mem\[2\]\[10\] _06566_ sky130_fd_sc_hd__mux2_2
X_21111_ VGND VPWR VPWR VGND _06007_ _02861_ keymem.key_mem\[6\]\[31\] _06008_ sky130_fd_sc_hd__mux2_2
XFILLER_0_67_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22091_ VGND VPWR _01758_ _06528_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21042_ VGND VPWR _05970_ _05969_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_5_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_10_584 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_242_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24801_ VGND VPWR VPWR VGND clk _01294_ reset_n keymem.key_mem\[6\]\[26\] sky130_fd_sc_hd__dfrtp_2
X_25781_ keymem.prev_key1_reg\[97\] clk _02274_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_242_947 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22993_ VGND VPWR VGND VPWR _02225_ _06963_ _06954_ keymem.prev_key1_reg\[48\] sky130_fd_sc_hd__o21a_2
XFILLER_0_173_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24732_ VGND VPWR VPWR VGND clk _01225_ reset_n keymem.key_mem\[7\]\[85\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_96_304 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21944_ VPWR VGND keymem.key_mem\[3\]\[37\] _06451_ _06439_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_171_1240 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_222_682 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24663_ VGND VPWR VPWR VGND clk _01156_ reset_n keymem.key_mem\[7\]\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_1029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21875_ VGND VPWR _06413_ _06405_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23614_ VGND VPWR VPWR VGND clk _00115_ reset_n keymem.key_mem\[14\]\[103\] sky130_fd_sc_hd__dfrtp_2
X_20826_ VGND VPWR VGND VPWR _05855_ keymem.key_mem_we _02743_ _05850_ _01166_ sky130_fd_sc_hd__a31o_2
XFILLER_0_166_236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24594_ VGND VPWR VPWR VGND clk _01087_ reset_n keymem.key_mem\[8\]\[75\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_437 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23545_ VGND VPWR VPWR VGND clk _00046_ reset_n keymem.key_mem\[14\]\[34\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20757_ VGND VPWR _01137_ _05815_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_110_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_174_280 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_24_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23476_ _07337_ _07339_ _03981_ _07338_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_107_347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20688_ VGND VPWR _01104_ _05779_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_169_1180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_64_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_122_1_Left_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25215_ VGND VPWR VPWR VGND clk _01708_ reset_n keymem.key_mem\[3\]\[56\] sky130_fd_sc_hd__dfrtp_2
X_22427_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[7\] _06707_ _06706_ _04889_ _01915_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_33_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13160_ VPWR VGND VPWR VGND keymem.key_mem\[4\]\[99\] _07734_ keymem.key_mem\[1\]\[99\]
+ _07558_ _08664_ sky130_fd_sc_hd__a22o_2
X_25146_ VGND VPWR VPWR VGND clk _01639_ reset_n keymem.key_mem\[4\]\[115\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_260_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22358_ VGND VPWR VPWR VGND _06669_ _03518_ keymem.key_mem\[2\]\[104\] _06670_ sky130_fd_sc_hd__mux2_2
XFILLER_0_108_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12111_ VGND VPWR VGND VPWR _07709_ _07580_ keymem.key_mem\[12\]\[5\] _07704_ _07708_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_260_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13091_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[92\] _07674_ keymem.key_mem\[1\]\[92\]
+ _07670_ _08602_ sky130_fd_sc_hd__a22o_2
X_21309_ VGND VPWR VPWR VGND _05971_ _03661_ keymem.key_mem\[6\]\[126\] _06111_ sky130_fd_sc_hd__mux2_2
XFILLER_0_130_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25077_ VGND VPWR VPWR VGND clk _01570_ reset_n keymem.key_mem\[4\]\[46\] sky130_fd_sc_hd__dfrtp_2
X_22289_ VGND VPWR _01851_ _06633_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12042_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[2\] _07535_ _07642_ _07635_ _07643_
+ sky130_fd_sc_hd__o22a_2
X_24028_ VGND VPWR VPWR VGND clk _00521_ reset_n keymem.key_mem\[12\]\[21\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_184_1_Left_451 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_79_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16850_ VGND VPWR VPWR VGND _02990_ _10963_ _02988_ _02691_ _02989_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_46_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_152_2_Left_623 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15801_ VGND VPWR _11257_ _11256_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16781_ VGND VPWR _02927_ _08936_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_219_1446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13993_ _09370_ _09465_ _09463_ _09464_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_219_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18520_ VGND VPWR VGND VPWR _04398_ _03951_ _04399_ _00316_ sky130_fd_sc_hd__a21o_2
X_15732_ enc_block.sword_ctr_reg\[1\] _11188_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[22\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_217_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12944_ VPWR VGND VPWR VGND _08468_ keymem.key_mem\[12\]\[78\] _07580_ keymem.key_mem\[4\]\[78\]
+ _07665_ _08469_ sky130_fd_sc_hd__a221o_2
XFILLER_0_137_1157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_220_619 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_217_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18451_ VPWR VGND VPWR VGND _04336_ block[66] _04330_ enc_block.block_w0_reg\[2\]
+ _04276_ _04337_ sky130_fd_sc_hd__a221o_2
XFILLER_0_73_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_87_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15663_ VPWR VGND VPWR VGND _11115_ _11119_ _11116_ _10673_ _11120_ sky130_fd_sc_hd__or4_2
XFILLER_0_241_991 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_213_1012 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_38_Left_306 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12875_ VPWR VGND VPWR VGND _08406_ keymem.key_mem\[14\]\[71\] _07782_ keymem.key_mem\[4\]\[71\]
+ _07914_ _08407_ sky130_fd_sc_hd__a221o_2
XFILLER_0_73_1189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17402_ VGND VPWR _00111_ _03486_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_157_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14614_ VGND VPWR VGND VPWR _10081_ _10080_ _10082_ keymem.prev_key0_reg\[4\] sky130_fd_sc_hd__a21oi_2
XFILLER_0_16_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11826_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[16\] dec_new_block\[80\]
+ _07477_ sky130_fd_sc_hd__mux2_2
X_18382_ VPWR VGND VPWR VGND _04275_ _04189_ _04273_ enc_block.block_w0_reg\[28\]
+ _03993_ _00302_ sky130_fd_sc_hd__a221o_2
X_15594_ VGND VPWR VPWR VGND _10378_ _11049_ key[142] _11052_ sky130_fd_sc_hd__mux2_2
XFILLER_0_200_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_258 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_95_381 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17333_ VPWR VGND VPWR VGND _03425_ _02677_ _03422_ key[219] _10838_ _03426_ sky130_fd_sc_hd__a221o_2
XFILLER_0_28_448 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14545_ VPWR VGND VPWR VGND _09150_ _10013_ _09656_ _09695_ sky130_fd_sc_hd__or3b_2
XFILLER_0_172_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11757_ VGND VPWR result[45] _07442_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_56_779 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17264_ VPWR VGND VPWR VGND _03363_ _10902_ _03361_ key[212] _03027_ _03364_ sky130_fd_sc_hd__a221o_2
XFILLER_0_102_12 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14476_ VGND VPWR VGND VPWR _09945_ _09005_ _09045_ _09044_ _09043_ sky130_fd_sc_hd__and4_2
X_11688_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[11\] dec_new_block\[11\]
+ _07408_ sky130_fd_sc_hd__mux2_2
X_19003_ VPWR VGND VPWR VGND _04832_ _04505_ enc_block.block_w2_reg\[26\] _04504_
+ _04833_ sky130_fd_sc_hd__a22o_2
X_16215_ VGND VPWR VGND VPWR _11270_ _11380_ _11464_ _02380_ sky130_fd_sc_hd__a21o_2
XFILLER_0_24_621 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13427_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[126\] _07872_ keymem.key_mem\[4\]\[126\]
+ _07636_ _08904_ sky130_fd_sc_hd__a22o_2
XFILLER_0_10_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17195_ VGND VPWR _03302_ _09512_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_125_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_148_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_440 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16146_ VGND VPWR VGND VPWR _11432_ _11596_ _11597_ _11598_ _11600_ _11599_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_84_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13358_ VPWR VGND VPWR VGND _08841_ keymem.key_mem\[5\]\[119\] _07683_ keymem.key_mem\[9\]\[119\]
+ _07738_ _08842_ sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_47_Left_315 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_267_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12309_ VGND VPWR _07893_ _07534_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16077_ VGND VPWR VGND VPWR _11520_ _11531_ _11532_ _11511_ _11526_ sky130_fd_sc_hd__nor4_2
X_13289_ VGND VPWR VGND VPWR _07841_ keymem.key_mem\[4\]\[112\] _08777_ _08779_ _08780_
+ _08736_ sky130_fd_sc_hd__a2111o_2
X_15028_ _10489_ _10492_ _10487_ _10491_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_19905_ VGND VPWR _00736_ _05364_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_18_Right_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_2_Left_555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_208_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19836_ VGND VPWR _05328_ _05246_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_237_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_999 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_120_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1018 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19767_ VGND VPWR _05292_ _05246_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16979_ VPWR VGND VPWR VGND _03107_ _02708_ _03104_ _03105_ _03106_ _10096_ sky130_fd_sc_hd__o311a_2
XFILLER_0_155_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18718_ VGND VPWR _04576_ _03957_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_127_86 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Left_324 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_91_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19698_ VGND VPWR VPWR VGND _05247_ keymem.key_mem\[11\]\[10\] _10836_ _05256_ sky130_fd_sc_hd__mux2_2
XFILLER_0_210_107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1279 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_56_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18649_ VGND VPWR _04515_ enc_block.block_w0_reg\[6\] _04514_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_1141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_78_359 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_91_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_318 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21660_ VGND VPWR _01557_ _06298_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_8_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_437 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20611_ VGND VPWR _01067_ _05739_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21591_ VGND VPWR _01525_ _06261_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_35_919 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23330_ VPWR VGND _07209_ _07208_ enc_block.round_key\[12\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_20542_ VGND VPWR _05703_ _05679_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_46_278 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_342 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23261_ VPWR VGND VGND VPWR _07126_ _07147_ _04042_ sky130_fd_sc_hd__nor2_2
X_20473_ VGND VPWR VPWR VGND _05660_ _03613_ keymem.key_mem\[9\]\[119\] _05666_ sky130_fd_sc_hd__mux2_2
XFILLER_0_229_1085 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25000_ VGND VPWR VPWR VGND clk _01493_ reset_n keymem.key_mem\[5\]\[97\] sky130_fd_sc_hd__dfrtp_2
X_22212_ VGND VPWR _01814_ _06593_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23192_ VGND VPWR VGND VPWR _07084_ _03664_ _03663_ _03667_ _07011_ sky130_fd_sc_hd__a211o_2
XFILLER_0_162_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_495 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22143_ VGND VPWR VPWR VGND _06554_ _09861_ keymem.key_mem\[2\]\[2\] _06557_ sky130_fd_sc_hd__mux2_2
XFILLER_0_24_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_203_1214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_190_2_Right_262 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Right_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22074_ VGND VPWR _01750_ _06519_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_168_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21025_ VGND VPWR VPWR VGND _05956_ _05075_ keymem.key_mem\[7\]\[120\] _05961_ sky130_fd_sc_hd__mux2_2
XFILLER_0_227_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25833_ VGND VPWR VPWR VGND clk _02326_ reset_n enc_block.block_w3_reg\[21\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_96_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_254_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_114 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25764_ keymem.prev_key1_reg\[80\] clk _02257_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22976_ VGND VPWR VGND VPWR _06953_ _02967_ _02966_ _02971_ _06951_ sky130_fd_sc_hd__a211o_2
XFILLER_0_74_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_134_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24715_ VGND VPWR VPWR VGND clk _01208_ reset_n keymem.key_mem\[7\]\[68\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_173_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21927_ VGND VPWR VGND VPWR _06441_ keymem.key_mem_we _02812_ _06432_ _01681_ sky130_fd_sc_hd__a31o_2
X_25695_ keymem.prev_key1_reg\[11\] clk _02188_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_179_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_74_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12660_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[50\] _07812_ keymem.key_mem\[11\]\[50\]
+ _07658_ _08213_ sky130_fd_sc_hd__a22o_2
X_24646_ VGND VPWR VPWR VGND clk _01139_ reset_n keymem.key_mem\[8\]\[127\] sky130_fd_sc_hd__dfrtp_2
X_21858_ VGND VPWR _06402_ _06401_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_33_1140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20809_ VGND VPWR VGND VPWR _05846_ keymem.key_mem_we _02340_ _05838_ _01158_ sky130_fd_sc_hd__a31o_2
X_12591_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[43\] _07748_ keymem.key_mem\[9\]\[43\]
+ _07672_ _08151_ sky130_fd_sc_hd__a22o_2
X_24577_ VGND VPWR VPWR VGND clk _01070_ reset_n keymem.key_mem\[8\]\[58\] sky130_fd_sc_hd__dfrtp_2
X_21789_ VGND VPWR _01619_ _06365_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_53_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14330_ VPWR VGND VPWR VGND _09800_ _09124_ sky130_fd_sc_hd__inv_2
X_23528_ VGND VPWR VPWR VGND clk _00029_ reset_n keymem.key_mem\[14\]\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_1425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_110_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14261_ VGND VPWR VPWR VGND _09730_ _09727_ key[130] _09731_ sky130_fd_sc_hd__mux2_2
XFILLER_0_0_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23459_ VPWR VGND VPWR VGND _07323_ block[26] _04139_ enc_block.block_w3_reg\[26\]
+ _04138_ _07324_ sky130_fd_sc_hd__a221o_2
XFILLER_0_11_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16000_ VGND VPWR _11455_ _11453_ _11454_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_184_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13212_ VPWR VGND VPWR VGND _08710_ keymem.key_mem\[3\]\[104\] _07619_ keymem.key_mem\[11\]\[104\]
+ _07838_ _08711_ sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_208_Left_475 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_81_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14192_ VPWR VGND VGND VPWR _09103_ _09663_ _09053_ sky130_fd_sc_hd__nor2_2
XFILLER_0_85_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_145_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_249_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_81_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25129_ VGND VPWR VPWR VGND clk _01622_ reset_n keymem.key_mem\[4\]\[98\] sky130_fd_sc_hd__dfrtp_2
X_13143_ VGND VPWR VGND VPWR _08649_ _08150_ keymem.key_mem\[3\]\[97\] _08646_ _08648_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_42_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_103_383 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_260_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_376 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17951_ VGND VPWR VPWR VGND _03896_ _03898_ keymem.prev_key0_reg\[107\] _03899_ sky130_fd_sc_hd__mux2_2
XFILLER_0_104_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13074_ VGND VPWR enc_block.round_key\[90\] _08586_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_221_1358 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_57_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16902_ VGND VPWR VGND VPWR _11539_ _11538_ _10386_ _03037_ sky130_fd_sc_hd__a21o_2
X_12025_ VGND VPWR VGND VPWR _07627_ _07619_ keymem.key_mem\[3\]\[1\] _07623_ _07626_
+ sky130_fd_sc_hd__a211o_2
X_17882_ VGND VPWR _00226_ _03851_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_206_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19621_ VGND VPWR _00603_ _05213_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_228_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_178_1279 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16833_ VGND VPWR VGND VPWR _10895_ _10894_ _02974_ _10896_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_258_1270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_195_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_73_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_217_Left_484 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19552_ VGND VPWR _00570_ _05177_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_191_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16764_ VGND VPWR VGND VPWR _02909_ _10088_ _02910_ _02911_ _02912_ keylen sky130_fd_sc_hd__a221oi_2
XFILLER_0_156_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13976_ VPWR VGND VGND VPWR _09416_ _09448_ _09380_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_63_Right_63 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_92_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_416 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_152_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15715_ VPWR VGND VPWR VGND _11171_ enc_block.block_w0_reg\[19\] _08951_ sky130_fd_sc_hd__or2_2
X_18503_ VPWR VGND _04384_ enc_block.block_w1_reg\[31\] enc_block.block_w1_reg\[30\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_53_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_191_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12927_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[76\] _07924_ keymem.key_mem\[4\]\[76\]
+ _08077_ _08454_ sky130_fd_sc_hd__a22o_2
XFILLER_0_232_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19483_ VGND VPWR VPWR VGND _05138_ _04931_ keymem.key_mem\[12\]\[38\] _05141_ sky130_fd_sc_hd__mux2_2
X_16695_ VGND VPWR _02848_ keymem.prev_key0_reg\[63\] keymem.prev_key0_reg\[95\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18434_ VGND VPWR _04321_ enc_block.block_w3_reg\[9\] _04320_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15646_ VGND VPWR VPWR VGND _09730_ _11101_ key[143] _11103_ sky130_fd_sc_hd__mux2_2
XFILLER_0_232_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12858_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[69\] _08391_ keymem.key_mem\[12\]\[69\]
+ _07673_ _08392_ sky130_fd_sc_hd__a22o_2
XFILLER_0_28_212 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11809_ VGND VPWR result[71] _07468_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18365_ VGND VPWR _04260_ _04259_ _04193_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15577_ VPWR VGND VGND VPWR _11036_ key[141] _10278_ sky130_fd_sc_hd__nand2_2
X_12789_ VPWR VGND VPWR VGND _08329_ keymem.key_mem\[6\]\[62\] _07711_ keymem.key_mem\[10\]\[62\]
+ _07785_ _08330_ sky130_fd_sc_hd__a221o_2
XFILLER_0_7_139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17316_ VGND VPWR _00101_ _03410_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_22_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14528_ VPWR VGND VPWR VGND _09994_ _09995_ _09996_ _09652_ _09964_ sky130_fd_sc_hd__or4b_2
XFILLER_0_125_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18296_ VGND VPWR VGND VPWR _04197_ _04196_ _04198_ _03966_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_113_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17247_ VGND VPWR _00094_ _03348_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_226_Left_493 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14459_ VGND VPWR VPWR VGND _09925_ keymem.prev_key1_reg\[67\] _09928_ _09927_ _09926_
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_163_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17178_ VGND VPWR _03287_ _03286_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_163_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_113_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_243_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16129_ VGND VPWR VGND VPWR _11578_ _11583_ _11580_ _11582_ _11579_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_60_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_690 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_209_774 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_209_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1368 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_100_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19819_ VGND VPWR _00695_ _05319_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22830_ VPWR VGND VPWR VGND _06862_ _08921_ _06861_ sky130_fd_sc_hd__or2_2
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_980 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_170_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_250_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22761_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[76\] _06837_ _06836_ _04992_ _02112_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24500_ VGND VPWR VPWR VGND clk _00993_ reset_n keymem.key_mem\[9\]\[109\] sky130_fd_sc_hd__dfrtp_2
X_21712_ VGND VPWR _01582_ _06325_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_211_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_250_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25480_ VGND VPWR VPWR VGND clk _01973_ reset_n keymem.key_mem\[1\]\[65\] sky130_fd_sc_hd__dfrtp_2
X_22692_ VGND VPWR VPWR VGND _06809_ keymem.key_mem\[0\]\[35\] _02904_ _06817_ sky130_fd_sc_hd__mux2_2
XFILLER_0_211_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24431_ VGND VPWR VPWR VGND clk _00924_ reset_n keymem.key_mem\[9\]\[40\] sky130_fd_sc_hd__dfrtp_2
X_21643_ VGND VPWR _01549_ _06289_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_170_50 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_351 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_110_1_Right_711 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24362_ VGND VPWR VPWR VGND clk _00855_ reset_n keymem.key_mem\[10\]\[99\] sky130_fd_sc_hd__dfrtp_2
X_21574_ VGND VPWR _01518_ _06251_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_191_367 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23313_ VPWR VGND VPWR VGND _07193_ _04874_ _07191_ enc_block.block_w3_reg\[10\]
+ _07115_ _02315_ sky130_fd_sc_hd__a221o_2
XFILLER_0_62_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20525_ VGND VPWR _01026_ _05694_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24293_ VGND VPWR VPWR VGND clk _00786_ reset_n keymem.key_mem\[10\]\[30\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_209_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_695 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_974 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23244_ VGND VPWR _07131_ enc_block.block_w3_reg\[28\] enc_block.block_w0_reg\[20\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20456_ VGND VPWR VPWR VGND _05649_ _03560_ keymem.key_mem\[9\]\[111\] _05657_ sky130_fd_sc_hd__mux2_2
XFILLER_0_127_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_203_1000 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_179_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20387_ VGND VPWR VPWR VGND _05614_ _03314_ keymem.key_mem\[9\]\[78\] _05621_ sky130_fd_sc_hd__mux2_2
X_23175_ VGND VPWR _02297_ _07073_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_28_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22126_ VGND VPWR _01775_ _06546_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_191_2_Right_263 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_184 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_219_538 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_98_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22057_ VGND VPWR VGND VPWR _06510_ keymem.key_mem_we _03418_ _06498_ _01742_ sky130_fd_sc_hd__a31o_2
XFILLER_0_265_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21008_ VGND VPWR VPWR VGND _05945_ _05058_ keymem.key_mem\[7\]\[112\] _05952_ sky130_fd_sc_hd__mux2_2
X_13830_ VGND VPWR _09302_ _09301_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25816_ VGND VPWR VPWR VGND clk _02309_ reset_n enc_block.block_w3_reg\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_138_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13761_ VPWR VGND VPWR VGND _09229_ _09063_ _09231_ _09232_ _09233_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_74_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25747_ keymem.prev_key1_reg\[63\] clk _02240_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_35_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22959_ VGND VPWR VPWR VGND _06914_ _06942_ keymem.prev_key1_reg\[35\] _06943_ sky130_fd_sc_hd__mux2_2
XFILLER_0_39_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15500_ VGND VPWR VGND VPWR _10533_ _10952_ _10956_ _10960_ _10959_ sky130_fd_sc_hd__nor4b_2
X_12712_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[55\] _08137_ keymem.key_mem\[11\]\[55\]
+ _07809_ _08260_ sky130_fd_sc_hd__a22o_2
XFILLER_0_74_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16480_ VGND VPWR VPWR VGND _02610_ _02638_ _02639_ _02641_ sky130_fd_sc_hd__or3_2
XFILLER_0_35_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13692_ VGND VPWR VGND VPWR _09164_ _09163_ _09152_ _09143_ _09131_ sky130_fd_sc_hd__and4_2
X_25678_ VGND VPWR VPWR VGND clk _02171_ reset_n keymem.rcon_logic.tmp_rcon\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_116_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_521 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15431_ VGND VPWR VGND VPWR _10874_ _10891_ _10892_ _10772_ _10881_ sky130_fd_sc_hd__nor4_2
XFILLER_0_2_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12643_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[48\] _07568_ keymem.key_mem\[2\]\[48\]
+ _07732_ _08198_ sky130_fd_sc_hd__a22o_2
XFILLER_0_210_1037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24629_ VGND VPWR VPWR VGND clk _01122_ reset_n keymem.key_mem\[8\]\[110\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_249_1225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_182_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_183 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_65_362 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18150_ VGND VPWR _04064_ _03955_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15362_ VGND VPWR VPWR VGND _10824_ _10823_ _10820_ _10821_ _09988_ sky130_fd_sc_hd__o31a_2
X_12574_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[42\] _07730_ keymem.key_mem\[12\]\[42\]
+ _07894_ _08135_ sky130_fd_sc_hd__a22o_2
X_17101_ VGND VPWR VPWR VGND _03185_ keymem.key_mem\[14\]\[67\] _03217_ _03218_ sky130_fd_sc_hd__mux2_2
XFILLER_0_0_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14313_ VGND VPWR _09782_ _09341_ _09783_ _09404_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_110_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_250 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_248 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18081_ _03999_ _04001_ _03982_ _04000_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_15293_ VPWR VGND VGND VPWR _10752_ _10753_ _10754_ _10755_ sky130_fd_sc_hd__nor3_2
XFILLER_0_29_1017 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_80_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_207 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17032_ VGND VPWR VPWR VGND _03153_ _02691_ _03155_ _09514_ _03154_ sky130_fd_sc_hd__o211a_2
XFILLER_0_145_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14244_ VPWR VGND VPWR VGND _09715_ keymem.prev_key0_reg\[1\] sky130_fd_sc_hd__inv_2
XFILLER_0_81_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_85_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14175_ VGND VPWR _09646_ _09166_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_1_849 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_81_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_46_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13126_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[96\] _07597_ keymem.key_mem\[3\]\[96\]
+ _08216_ _08633_ sky130_fd_sc_hd__a22o_2
XFILLER_0_239_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18983_ VGND VPWR _04815_ enc_block.block_w1_reg\[0\] _04753_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_264_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17934_ VGND VPWR VPWR VGND _03876_ key[230] keymem.prev_key1_reg\[102\] _03887_
+ sky130_fd_sc_hd__mux2_2
X_13057_ VGND VPWR VGND VPWR _07780_ keymem.key_mem\[5\]\[89\] _08568_ _08570_ _08571_
+ _08480_ sky130_fd_sc_hd__a2111o_2
XPHY_EDGE_ROW_65_2_Right_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12008_ VGND VPWR _07610_ _07609_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_84_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_733 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17865_ VGND VPWR VPWR VGND _03812_ key[208] keymem.prev_key1_reg\[80\] _03840_ sky130_fd_sc_hd__mux2_2
X_19604_ VGND VPWR VGND VPWR _05204_ keymem.key_mem_we _03460_ _05187_ _00595_ sky130_fd_sc_hd__a31o_2
X_16816_ VPWR VGND VPWR VGND _02959_ key[41] _09987_ sky130_fd_sc_hd__or2_2
XFILLER_0_117_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_191_1232 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_147_1_Left_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17796_ VGND VPWR _03793_ _02947_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_156_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19535_ VGND VPWR VGND VPWR _05168_ keymem.key_mem_we _03173_ _05164_ _00562_ sky130_fd_sc_hd__a31o_2
X_13959_ VGND VPWR _09431_ _09430_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_92_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16747_ VGND VPWR VPWR VGND _10091_ key[163] keymem.prev_key1_reg\[35\] _02896_ sky130_fd_sc_hd__mux2_2
XFILLER_0_117_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19466_ VGND VPWR VGND VPWR _05131_ keymem.key_mem_we _02839_ _05121_ _00530_ sky130_fd_sc_hd__a31o_2
X_16678_ VGND VPWR VGND VPWR _02829_ _02830_ _02832_ _02828_ sky130_fd_sc_hd__nand3_2
XFILLER_0_18_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18417_ VPWR VGND VGND VPWR _04305_ _04304_ enc_block.sword_ctr_reg\[1\] _08923_
+ _07394_ _00307_ sky130_fd_sc_hd__a311o_2
XFILLER_0_232_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15629_ VGND VPWR VPWR VGND _11086_ _11087_ _11085_ _11081_ _10668_ _10593_ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_158_386 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19397_ VGND VPWR _05093_ _05092_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_5_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_234_Left_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18348_ VGND VPWR VGND VPWR _04244_ _04243_ _04245_ _03966_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_16_226 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_267_1369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18279_ VGND VPWR _04182_ _04110_ _04181_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_44_579 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20310_ VGND VPWR VPWR VGND _05580_ _02964_ keymem.key_mem\[9\]\[41\] _05581_ sky130_fd_sc_hd__mux2_2
XFILLER_0_128_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_163_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21290_ VGND VPWR _01384_ _06101_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_3_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_124_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20241_ VGND VPWR _00892_ _05544_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_163_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1391 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_64_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20172_ VGND VPWR _00861_ _05506_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_99_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_255_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_243_Left_510 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_196_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24980_ VGND VPWR VPWR VGND clk _01473_ reset_n keymem.key_mem\[5\]\[77\] sky130_fd_sc_hd__dfrtp_2
X_23931_ VGND VPWR VPWR VGND clk _00424_ reset_n keymem.key_mem\[13\]\[52\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_239_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_79_1_Left_346 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_100_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_552 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23862_ VGND VPWR VPWR VGND clk _00355_ reset_n enc_block.block_w2_reg\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_224_563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_131_1_Left_398 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_174_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25601_ VGND VPWR VPWR VGND clk _02094_ reset_n keymem.key_mem\[0\]\[58\] sky130_fd_sc_hd__dfrtp_2
X_22813_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[112\] _06860_ _06859_ _05058_ _02148_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_196_415 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23793_ VGND VPWR VPWR VGND clk _00286_ reset_n enc_block.block_w0_reg\[12\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_75_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25532_ VGND VPWR VPWR VGND clk _02025_ reset_n keymem.key_mem\[1\]\[117\] sky130_fd_sc_hd__dfrtp_2
X_22744_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[66\] _06837_ _06836_ _04977_ _02102_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_39_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_0_Right_0 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_215_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25463_ VGND VPWR VPWR VGND clk _01956_ reset_n keymem.key_mem\[1\]\[48\] sky130_fd_sc_hd__dfrtp_2
X_22675_ VGND VPWR _06809_ _06784_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_133_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_211_1368 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_109_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24414_ VGND VPWR VPWR VGND clk _00907_ reset_n keymem.key_mem\[9\]\[23\] sky130_fd_sc_hd__dfrtp_2
X_21626_ VGND VPWR _01541_ _06280_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_164_345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_63_833 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_193_1_Left_460 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25394_ VGND VPWR VPWR VGND clk _01887_ reset_n keymem.key_mem\[2\]\[107\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_535 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_62_321 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_124_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_332 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_8_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_1_Right_712 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_111_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24345_ VGND VPWR VPWR VGND clk _00838_ reset_n keymem.key_mem\[10\]\[82\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_161_2_Left_632 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21557_ VGND VPWR VPWR VGND _06242_ _03580_ keymem.key_mem\[5\]\[114\] _06243_ sky130_fd_sc_hd__mux2_2
XFILLER_0_62_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20508_ VGND VPWR _01018_ _05685_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_181_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12290_ VGND VPWR _07876_ _07674_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24276_ VGND VPWR VPWR VGND clk _00769_ reset_n keymem.key_mem\[10\]\[13\] sky130_fd_sc_hd__dfrtp_2
X_21488_ VGND VPWR _01477_ _06206_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_15_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_590 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_741 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_107_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_142_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23227_ VGND VPWR _07115_ _07093_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20439_ VGND VPWR VPWR VGND _05638_ _03511_ keymem.key_mem\[9\]\[103\] _05648_ sky130_fd_sc_hd__mux2_2
XFILLER_0_200_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_31_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23158_ VGND VPWR _02290_ _07063_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_222_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22109_ VGND VPWR _01767_ _06537_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_192_2_Right_264 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15980_ VPWR VGND VPWR VGND _11435_ _11433_ _11407_ _11409_ _11432_ _11436_ sky130_fd_sc_hd__a221o_2
XFILLER_0_257_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23089_ VGND VPWR VGND VPWR _07020_ _03398_ _06891_ _03400_ _07011_ sky130_fd_sc_hd__a211o_2
XFILLER_0_179_1363 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_1148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14931_ VGND VPWR VGND VPWR enc_block.block_w1_reg\[8\] _08947_ _10387_ _10393_ _10395_
+ _10394_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_257_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_861 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14862_ VGND VPWR _10327_ _08936_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17650_ VGND VPWR VPWR VGND _03691_ key[137] keymem.prev_key1_reg\[9\] _03696_ sky130_fd_sc_hd__mux2_2
XFILLER_0_54_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13813_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[29\] _08969_ _09285_ _08964_ _09283_
+ _09284_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_216_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16601_ VGND VPWR VGND VPWR _02756_ keymem.prev_key1_reg\[91\] _02758_ _02755_ sky130_fd_sc_hd__nand3_2
XFILLER_0_230_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17581_ VGND VPWR _00135_ _03641_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14793_ _10257_ _10259_ _10256_ _10258_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_225_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_153_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16532_ VGND VPWR _02691_ _09717_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19320_ VGND VPWR _00475_ _05040_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13744_ VGND VPWR _09216_ _09210_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_11_Left_279 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_1054 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16463_ VGND VPWR VGND VPWR _11270_ _11308_ _11267_ _11330_ _02624_ sky130_fd_sc_hd__o22a_2
XFILLER_0_6_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19251_ VPWR VGND keymem.key_mem_we _04997_ _03314_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13675_ VPWR VGND VPWR VGND _09044_ _09005_ _09034_ _09001_ _09147_ sky130_fd_sc_hd__or4_2
XFILLER_0_2_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15414_ VPWR VGND VGND VPWR _10602_ _10875_ _10520_ sky130_fd_sc_hd__nor2_2
X_18202_ VGND VPWR _04112_ _04109_ _04111_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_513 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12626_ VGND VPWR enc_block.round_key\[46\] _08182_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19182_ VGND VPWR VPWR VGND _04951_ _04955_ keymem.key_mem\[13\]\[50\] _04956_ sky130_fd_sc_hd__mux2_2
XFILLER_0_155_345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16394_ VPWR VGND VPWR VGND _02554_ _02555_ _02556_ _11568_ _02553_ sky130_fd_sc_hd__or4b_2
XPHY_EDGE_ROW_93_2_Left_564 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_264_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_155_378 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18133_ _04047_ _04049_ _04008_ _04048_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_15345_ VGND VPWR VGND VPWR _10611_ _10507_ _10807_ _10602_ sky130_fd_sc_hd__a21oi_2
X_12557_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[40\] _08096_ keymem.key_mem\[12\]\[40\]
+ _07808_ _08120_ sky130_fd_sc_hd__a22o_2
XFILLER_0_79_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18064_ VPWR VGND _03985_ enc_block.block_w0_reg\[25\] enc_block.block_w1_reg\[17\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_227_1353 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15276_ VGND VPWR keymem.prev_key1_reg\[73\] _10737_ _10739_ _10738_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_12488_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[34\] _07650_ keymem.key_mem\[12\]\[34\]
+ _07788_ _08057_ sky130_fd_sc_hd__a22o_2
XFILLER_0_41_549 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17015_ VGND VPWR _03140_ _03139_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_160_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14227_ VPWR VGND VGND VPWR _09216_ _09138_ _09698_ _09116_ _09122_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_21_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_288 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_46_1183 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14158_ VGND VPWR VGND VPWR _09598_ _09628_ _09629_ _09438_ _09606_ sky130_fd_sc_hd__nor4_2
XFILLER_0_240_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13109_ VGND VPWR VGND VPWR _08016_ keymem.key_mem\[7\]\[94\] _08615_ _08617_ _08618_
+ _08599_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_201_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14089_ VGND VPWR VPWR VGND _09468_ _09305_ _09559_ _09560_ sky130_fd_sc_hd__or3_2
X_18966_ VGND VPWR _04800_ enc_block.block_w0_reg\[14\] _04799_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_237_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17917_ VGND VPWR _00237_ _03875_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_66_2_Right_138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18897_ VPWR VGND VPWR VGND _04738_ _04736_ _04737_ sky130_fd_sc_hd__or2_2
XFILLER_0_28_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_861 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17848_ VGND VPWR _00215_ _03828_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_234_1313 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_156_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_221_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17779_ VGND VPWR VPWR VGND _03719_ key[181] keymem.prev_key1_reg\[53\] _03781_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19518_ VGND VPWR VGND VPWR _05159_ keymem.key_mem_we _03091_ _05135_ _00554_ sky130_fd_sc_hd__a31o_2
X_20790_ VPWR VGND keymem.key_mem\[7\]\[10\] _05836_ _05830_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_14_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19449_ VGND VPWR VGND VPWR _05122_ keymem.key_mem_we _02608_ _05121_ _00522_ sky130_fd_sc_hd__a31o_2
XFILLER_0_146_312 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_29_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22460_ VGND VPWR VPWR VGND _06715_ keymem.key_mem\[1\]\[24\] _02689_ _06724_ sky130_fd_sc_hd__mux2_2
XFILLER_0_9_779 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_88_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21411_ VGND VPWR _01440_ _06166_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_45_866 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_97_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22391_ VGND VPWR VPWR VGND _06680_ _03620_ keymem.key_mem\[2\]\[120\] _06687_ sky130_fd_sc_hd__mux2_2
XFILLER_0_267_1199 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_161_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24130_ VGND VPWR VPWR VGND clk _00623_ reset_n keymem.key_mem\[12\]\[123\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_440 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_527 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21342_ VGND VPWR _06130_ _10913_ _01407_ _06114_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_60_858 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_128_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24061_ VGND VPWR VPWR VGND clk _00554_ reset_n keymem.key_mem\[12\]\[54\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_495 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21273_ VGND VPWR _01376_ _06092_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_128_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23012_ VGND VPWR VPWR VGND _02233_ _03103_ _03107_ _06925_ _06974_ sky130_fd_sc_hd__o31a_2
XFILLER_0_60_1114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20224_ VGND VPWR VPWR VGND _05535_ _09537_ keymem.key_mem\[9\]\[0\] _05536_ sky130_fd_sc_hd__mux2_2
XFILLER_0_25_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_99_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20155_ VGND VPWR _00853_ _05497_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_25_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_99_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20086_ VGND VPWR _00820_ _05461_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24963_ VGND VPWR VPWR VGND clk _01456_ reset_n keymem.key_mem\[5\]\[60\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_1010 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23914_ VGND VPWR VPWR VGND clk _00407_ reset_n keymem.key_mem\[13\]\[35\] sky130_fd_sc_hd__dfrtp_2
X_24894_ VGND VPWR VPWR VGND clk _01387_ reset_n keymem.key_mem\[6\]\[119\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_135_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23845_ VGND VPWR VPWR VGND clk _00338_ reset_n enc_block.block_w1_reg\[30\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_139_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_746 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_197_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_135_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_566 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11790_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[30\] dec_new_block\[62\]
+ _07459_ sky130_fd_sc_hd__mux2_2
X_23776_ VGND VPWR VPWR VGND clk _00269_ reset_n enc_block.round\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_170_1157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20988_ VGND VPWR _01242_ _05941_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_32_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_36_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25515_ VGND VPWR VPWR VGND clk _02008_ reset_n keymem.key_mem\[1\]\[100\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_211_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22727_ VGND VPWR _02094_ _06828_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13460_ VPWR VGND _08932_ _08931_ keymem.prev_key0_reg\[0\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_25446_ VGND VPWR VPWR VGND clk _01939_ reset_n keymem.key_mem\[1\]\[31\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_94_298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22658_ VGND VPWR _02053_ _06800_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_63_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12411_ VPWR VGND VPWR VGND _07986_ keymem.key_mem\[6\]\[27\] _07565_ keymem.key_mem\[2\]\[27\]
+ _07646_ _07987_ sky130_fd_sc_hd__a221o_2
X_21609_ VGND VPWR _01533_ _06271_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25377_ VGND VPWR VPWR VGND clk _01870_ reset_n keymem.key_mem\[2\]\[90\] sky130_fd_sc_hd__dfrtp_2
X_13391_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[122\] _07612_ keymem.key_mem\[1\]\[122\]
+ _07670_ _08872_ sky130_fd_sc_hd__a22o_2
XFILLER_0_211_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22589_ VGND VPWR _06775_ _06696_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15130_ VPWR VGND VPWR VGND _10457_ _10435_ _10430_ _10443_ _10594_ sky130_fd_sc_hd__or4_2
XFILLER_0_50_302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_685 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_112_1_Right_713 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24328_ VGND VPWR VPWR VGND clk _00821_ reset_n keymem.key_mem\[10\]\[65\] sky130_fd_sc_hd__dfrtp_2
X_12342_ VGND VPWR _07924_ _07592_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_69_1194 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_146_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15061_ VPWR VGND VGND VPWR _10524_ _10525_ _10504_ sky130_fd_sc_hd__nor2_2
XFILLER_0_50_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24259_ VGND VPWR VPWR VGND clk _00752_ reset_n keymem.key_mem\[11\]\[124\] sky130_fd_sc_hd__dfrtp_2
X_12273_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[16\] _07592_ keymem.key_mem\[2\]\[16\]
+ _07732_ _07860_ sky130_fd_sc_hd__a22o_2
XFILLER_0_43_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14012_ VGND VPWR VGND VPWR _09426_ _09415_ _09386_ _09411_ _09484_ sky130_fd_sc_hd__o22a_2
XFILLER_0_47_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_931 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_107_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18820_ VGND VPWR _04669_ enc_block.block_w1_reg\[6\] _04668_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_193_2_Right_265 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18751_ VPWR VGND _04606_ enc_block.block_w2_reg\[25\] enc_block.block_w3_reg\[17\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_15963_ VPWR VGND VPWR VGND _11173_ _11221_ _11247_ _11166_ _11419_ sky130_fd_sc_hd__or4_2
XFILLER_0_65_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17702_ VGND VPWR _03733_ _03679_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14914_ VGND VPWR _10378_ _09729_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15894_ VPWR VGND VPWR VGND _11230_ _11349_ _11292_ _11348_ _11350_ sky130_fd_sc_hd__a22o_2
X_18682_ VGND VPWR _04544_ enc_block.block_w0_reg\[2\] _04331_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_17633_ VGND VPWR _00144_ _03684_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_118_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14845_ VGND VPWR VGND VPWR _09444_ _09564_ _09381_ _09749_ _10310_ sky130_fd_sc_hd__o22a_2
XFILLER_0_157_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_341 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_216_1065 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_54_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14776_ VPWR VGND VGND VPWR _09385_ _10237_ _10239_ _10241_ _10242_ sky130_fd_sc_hd__and4b_2
XFILLER_0_19_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17564_ VPWR VGND VPWR VGND _03626_ _03623_ _03622_ key[249] _08929_ _03627_ sky130_fd_sc_hd__a221o_2
X_11988_ VGND VPWR _07591_ _07590_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_114_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19303_ VPWR VGND keymem.key_mem_we _05029_ _03480_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_54_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13727_ VGND VPWR VGND VPWR _09199_ _09005_ _08991_ _09044_ _09043_ sky130_fd_sc_hd__and4_2
XFILLER_0_188_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16515_ VGND VPWR _02675_ _02672_ _02674_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_17495_ VPWR VGND VPWR VGND _03566_ _03494_ _03562_ key[240] _03527_ _03567_ sky130_fd_sc_hd__a221o_2
XFILLER_0_6_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19234_ VPWR VGND keymem.key_mem_we _04986_ _03259_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13658_ VGND VPWR VGND VPWR _09127_ _09128_ _09129_ _09125_ _09130_ sky130_fd_sc_hd__o22a_2
X_16446_ VGND VPWR _02608_ _02607_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_89_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_264_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12609_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[45\] _07984_ keymem.key_mem\[2\]\[45\]
+ _07547_ _08167_ sky130_fd_sc_hd__a22o_2
XFILLER_0_229_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16377_ VGND VPWR VPWR VGND keymem.prev_key0_reg\[117\] _02538_ _02540_ _02537_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_121_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19165_ VGND VPWR _00416_ _04944_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13589_ VGND VPWR VGND VPWR _09061_ _09015_ _09045_ _09014_ _09043_ sky130_fd_sc_hd__and4_2
XFILLER_0_87_1250 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_30_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15328_ VPWR VGND VPWR VGND _10790_ _10496_ _10527_ sky130_fd_sc_hd__or2_2
X_18116_ VPWR VGND _04033_ enc_block.block_w0_reg\[28\] enc_block.block_w3_reg\[4\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_205_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19096_ VGND VPWR VGND VPWR _04902_ keymem.key_mem_we _11547_ _04896_ _00389_ sky130_fd_sc_hd__a31o_2
XFILLER_0_129_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15259_ VPWR VGND VGND VPWR _10538_ _10722_ _10609_ sky130_fd_sc_hd__nor2_2
X_18047_ VPWR VGND _03969_ _03968_ enc_block.round_key\[96\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_125_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_205_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_777 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_22_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19998_ VGND VPWR _00778_ _05415_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_201_1345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_96_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18949_ VPWR VGND VGND VPWR _04784_ _04785_ _04382_ sky130_fd_sc_hd__nor2_2
XFILLER_0_254_967 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_214_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_197_1282 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_67_2_Right_139 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21960_ VGND VPWR VPWR VGND _06449_ _04945_ keymem.key_mem\[3\]\[45\] _06459_ sky130_fd_sc_hd__mux2_2
XFILLER_0_20_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_146_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20911_ VGND VPWR _01205_ _05901_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_146_96 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21891_ VPWR VGND keymem.key_mem\[3\]\[13\] _06422_ _06413_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_402 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23630_ VGND VPWR VPWR VGND clk _00131_ reset_n keymem.key_mem\[14\]\[119\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_136_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20842_ VGND VPWR _05864_ _05820_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_230_1018 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_162_40 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_221_396 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23561_ VGND VPWR VPWR VGND clk _00062_ reset_n keymem.key_mem\[14\]\[50\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_212_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20773_ VPWR VGND keymem.key_mem\[7\]\[2\] _05827_ _05824_ VPWR VGND sky130_fd_sc_hd__and2_2
X_25300_ VGND VPWR VPWR VGND clk _01793_ reset_n keymem.key_mem\[2\]\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_146_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22512_ VGND VPWR _01964_ _06743_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_71_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23492_ VPWR VGND VPWR VGND _07352_ _04065_ enc_block.block_w3_reg\[30\] _03953_
+ _07353_ sky130_fd_sc_hd__a22o_2
XFILLER_0_64_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25231_ VGND VPWR VPWR VGND clk _01724_ reset_n keymem.key_mem\[3\]\[72\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22443_ VGND VPWR _06715_ _06701_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_45_663 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_91_268 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_146_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_18_888 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_814 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25162_ VGND VPWR VPWR VGND clk _01655_ reset_n keymem.key_mem\[3\]\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_324 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22374_ VGND VPWR VPWR VGND _06669_ _03567_ keymem.key_mem\[2\]\[112\] _06678_ sky130_fd_sc_hd__mux2_2
X_24113_ VGND VPWR VPWR VGND clk _00606_ reset_n keymem.key_mem\[12\]\[106\] sky130_fd_sc_hd__dfrtp_2
X_21325_ VGND VPWR _01399_ _06121_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25093_ VGND VPWR VPWR VGND clk _01586_ reset_n keymem.key_mem\[4\]\[62\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_143_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_292 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24044_ VGND VPWR VPWR VGND clk _00537_ reset_n keymem.key_mem\[12\]\[37\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_104_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21256_ VGND VPWR _01368_ _06083_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_223_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20207_ VGND VPWR _00878_ _05524_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21187_ VGND VPWR _01335_ _06047_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_229_474 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_257_794 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20138_ VGND VPWR _00845_ _05488_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24946_ VGND VPWR VPWR VGND clk _01439_ reset_n keymem.key_mem\[5\]\[43\] sky130_fd_sc_hd__dfrtp_2
X_12960_ VPWR VGND VPWR VGND _08483_ keymem.key_mem\[13\]\[79\] _07730_ keymem.key_mem\[12\]\[79\]
+ _07894_ _08484_ sky130_fd_sc_hd__a221o_2
X_20069_ VGND VPWR _00812_ _05452_ VPWR VGND sky130_fd_sc_hd__buf_1
X_11911_ VGND VPWR result[122] _07519_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24877_ VGND VPWR VPWR VGND clk _01370_ reset_n keymem.key_mem\[6\]\[102\] sky130_fd_sc_hd__dfrtp_2
X_12891_ VGND VPWR enc_block.round_key\[72\] _08421_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14630_ VPWR VGND VPWR VGND _10097_ _10085_ _10084_ key[132] _09544_ _10098_ sky130_fd_sc_hd__a221o_2
X_23828_ VGND VPWR VPWR VGND clk _00321_ reset_n enc_block.block_w1_reg\[13\] sky130_fd_sc_hd__dfrtp_2
X_11842_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[24\] dec_new_block\[88\]
+ _07485_ sky130_fd_sc_hd__mux2_2
XFILLER_0_213_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_197_587 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14561_ VGND VPWR _10028_ _09168_ _10029_ _09160_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_32_1013 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23759_ keymem.prev_key0_reg\[115\] clk _00256_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_11773_ VGND VPWR result[53] _07450_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_230_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13512_ VPWR VGND VGND VPWR enc_block.block_w1_reg\[5\] enc_block.sword_ctr_reg\[0\]
+ _08984_ sky130_fd_sc_hd__or2b_2
X_16300_ VGND VPWR VGND VPWR _02462_ _02460_ _02464_ _02461_ sky130_fd_sc_hd__nand3_2
X_17280_ VGND VPWR VGND VPWR _03377_ _03376_ _10386_ _03378_ sky130_fd_sc_hd__a21o_2
X_14492_ VGND VPWR VGND VPWR _09961_ _09060_ _09184_ _09135_ sky130_fd_sc_hd__and3b_2
XFILLER_0_55_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_198_Right_67 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16231_ VGND VPWR _02396_ keymem.prev_key0_reg\[115\] _02395_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_13443_ VGND VPWR VGND VPWR _08919_ _07842_ keymem.key_mem\[9\]\[127\] _08916_ _08918_
+ sky130_fd_sc_hd__a211o_2
X_25429_ VGND VPWR VPWR VGND clk _01922_ reset_n keymem.key_mem\[1\]\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_125_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16162_ VGND VPWR VGND VPWR _11616_ _11407_ _11340_ _11348_ _11417_ _11396_ sky130_fd_sc_hd__a32o_2
XFILLER_0_207_1009 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13374_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[120\] _08027_ _08856_ _08852_ _08857_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_63_493 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_24_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15113_ VGND VPWR _10576_ _10455_ _10577_ _10572_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_113_1_Right_714 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12325_ VGND VPWR _07908_ _07771_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_156_1_Left_423 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16093_ VGND VPWR VPWR VGND _11041_ keymem.key_mem\[14\]\[17\] _11547_ _11548_ sky130_fd_sc_hd__mux2_2
X_15044_ VGND VPWR _10508_ _10507_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19921_ VGND VPWR VPWR VGND _05372_ keymem.key_mem\[11\]\[116\] _03592_ _05373_ sky130_fd_sc_hd__mux2_2
X_12256_ VGND VPWR _07845_ _07613_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_255_709 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19852_ VGND VPWR _00711_ _05336_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12187_ VGND VPWR _07780_ _07779_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18803_ VGND VPWR _04654_ _04599_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_247_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_78_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19783_ VGND VPWR _00678_ _05300_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_247_73 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16995_ VPWR VGND _03121_ _02729_ _02728_ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_120_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_223_606 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_207_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_194_2_Right_266 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18734_ VPWR VGND VPWR VGND _04590_ _04550_ _04589_ enc_block.block_w1_reg\[31\]
+ _04328_ _00339_ sky130_fd_sc_hd__a221o_2
X_15946_ VGND VPWR VGND VPWR _11402_ _11222_ _11395_ _11167_ _11266_ sky130_fd_sc_hd__a211o_2
XFILLER_0_92_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_28 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_820 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_216_691 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18665_ VPWR VGND _04529_ _04306_ enc_block.block_w1_reg\[31\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15877_ VPWR VGND VGND VPWR _11325_ _11327_ _11333_ _11332_ _11330_ sky130_fd_sc_hd__o22ai_2
X_17616_ VGND VPWR VGND VPWR _09524_ keymem.prev_key1_reg\[0\] _03671_ _03670_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_155_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14828_ VGND VPWR VGND VPWR _09399_ _09294_ _09475_ _09392_ _10293_ sky130_fd_sc_hd__o22a_2
X_18596_ VGND VPWR VGND VPWR _04467_ _04266_ _04316_ _04468_ enc_block.block_w1_reg\[16\]
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_118_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_19_608 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17547_ VPWR VGND _09533_ _03612_ _03611_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_15_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14759_ VGND VPWR VGND VPWR _09109_ _09136_ _10225_ _09067_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_188_1215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_89_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17478_ VGND VPWR VPWR VGND _11456_ _11047_ key[238] _03552_ sky130_fd_sc_hd__mux2_2
X_19217_ VGND VPWR VPWR VGND _04951_ _04975_ keymem.key_mem\[13\]\[65\] _04976_ sky130_fd_sc_hd__mux2_2
XFILLER_0_89_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16429_ VGND VPWR VGND VPWR _02590_ _02591_ _02589_ _02588_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_128_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_460 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_88_1_Left_355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_264_1158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19148_ VPWR VGND keymem.key_mem_we _04933_ _02945_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_30_806 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19079_ VPWR VGND keymem.key_mem\[13\]\[10\] _04893_ _04887_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_41_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21110_ VGND VPWR _06007_ _05971_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_1_240 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22090_ VGND VPWR VPWR VGND _06527_ _05045_ keymem.key_mem\[3\]\[106\] _06528_ sky130_fd_sc_hd__mux2_2
XFILLER_0_1_262 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_10_541 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_284 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_552 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21041_ VGND VPWR VGND VPWR _05969_ keymem.round_ctr_reg\[2\] _05385_ keymem.round_ctr_reg\[3\]
+ sky130_fd_sc_hd__and3b_2
XFILLER_0_201_1186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24800_ VGND VPWR VPWR VGND clk _01293_ reset_n keymem.key_mem\[6\]\[25\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_226_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25780_ keymem.prev_key1_reg\[96\] clk _02273_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22992_ VGND VPWR VGND VPWR _06963_ _03031_ _03028_ _03034_ _06951_ sky130_fd_sc_hd__a211o_2
XFILLER_0_198_318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24731_ VGND VPWR VPWR VGND clk _01224_ reset_n keymem.key_mem\[7\]\[84\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_170_2_Left_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21943_ VGND VPWR _01688_ _06450_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_171_1230 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24662_ VGND VPWR VPWR VGND clk _01155_ reset_n keymem.key_mem\[7\]\[15\] sky130_fd_sc_hd__dfrtp_2
X_21874_ VGND VPWR VGND VPWR _06412_ keymem.key_mem_we _10194_ _06404_ _01657_ sky130_fd_sc_hd__a31o_2
XFILLER_0_173_83 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_210_834 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23613_ VGND VPWR VPWR VGND clk _00114_ reset_n keymem.key_mem\[14\]\[102\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_210_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20825_ VPWR VGND keymem.key_mem\[7\]\[26\] _05855_ _05844_ VPWR VGND sky130_fd_sc_hd__and2_2
X_24593_ VGND VPWR VPWR VGND clk _01086_ reset_n keymem.key_mem\[8\]\[74\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_166_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_340 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23544_ VGND VPWR VPWR VGND clk _00045_ reset_n keymem.key_mem\[14\]\[33\] sky130_fd_sc_hd__dfrtp_2
X_20756_ VGND VPWR VPWR VGND _05805_ _03654_ keymem.key_mem\[8\]\[125\] _05815_ sky130_fd_sc_hd__mux2_2
XFILLER_0_37_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_68_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23475_ VPWR VGND VPWR VGND _07338_ _07130_ _07336_ sky130_fd_sc_hd__or2_2
XFILLER_0_107_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20687_ VGND VPWR VPWR VGND _05772_ _03434_ keymem.key_mem\[8\]\[92\] _05779_ sky130_fd_sc_hd__mux2_2
XFILLER_0_107_359 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25214_ VGND VPWR VPWR VGND clk _01707_ reset_n keymem.key_mem\[3\]\[55\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_220_Right_89 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22426_ VGND VPWR _06707_ _06696_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_32_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25145_ VGND VPWR VPWR VGND clk _01638_ reset_n keymem.key_mem\[4\]\[114\] sky130_fd_sc_hd__dfrtp_2
X_22357_ VGND VPWR _06669_ _06552_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_32_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12110_ VPWR VGND VPWR VGND _07707_ keymem.key_mem\[14\]\[5\] _07706_ keymem.key_mem\[9\]\[5\]
+ _07705_ _07708_ sky130_fd_sc_hd__a221o_2
XFILLER_0_108_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21308_ VGND VPWR _01393_ _06110_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_206_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13090_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[92\] _07725_ keymem.key_mem\[14\]\[92\]
+ _07666_ _08601_ sky130_fd_sc_hd__a22o_2
X_25076_ VGND VPWR VPWR VGND clk _01569_ reset_n keymem.key_mem\[4\]\[45\] sky130_fd_sc_hd__dfrtp_2
X_22288_ VGND VPWR VPWR VGND _06622_ _03251_ keymem.key_mem\[2\]\[71\] _06633_ sky130_fd_sc_hd__mux2_2
X_24027_ VGND VPWR VPWR VGND clk _00520_ reset_n keymem.key_mem\[12\]\[20\] sky130_fd_sc_hd__dfrtp_2
X_12041_ VGND VPWR VGND VPWR _07642_ _07610_ keymem.key_mem\[7\]\[2\] _07638_ _07641_
+ sky130_fd_sc_hd__a211o_2
X_21239_ VGND VPWR _01360_ _06074_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_79_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15800_ VPWR VGND VPWR VGND _11192_ _11208_ _11207_ _11187_ _11256_ sky130_fd_sc_hd__or4_2
XFILLER_0_260_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13992_ VGND VPWR VGND VPWR _09464_ _09291_ _09339_ _09328_ _09306_ sky130_fd_sc_hd__and4_2
X_16780_ VGND VPWR VGND VPWR _10267_ _10266_ _02691_ _02926_ sky130_fd_sc_hd__a21o_2
XFILLER_0_258_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15731_ VGND VPWR VGND VPWR _11187_ _11186_ _11185_ keymem.prev_key1_reg\[23\] _10402_
+ _09255_ sky130_fd_sc_hd__a32o_2
X_12943_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[78\] _07912_ keymem.key_mem\[10\]\[78\]
+ _07629_ _08468_ sky130_fd_sc_hd__a22o_2
XFILLER_0_176_1185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_1222 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24929_ VGND VPWR VPWR VGND clk _01422_ reset_n keymem.key_mem\[5\]\[26\] sky130_fd_sc_hd__dfrtp_2
X_18450_ _04334_ _04336_ _04294_ _04335_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_15662_ VGND VPWR VGND VPWR _11119_ _10515_ _10638_ _11117_ _11118_ sky130_fd_sc_hd__a211o_2
XFILLER_0_62_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12874_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[71\] _07918_ keymem.key_mem\[12\]\[71\]
+ _07806_ _08406_ sky130_fd_sc_hd__a22o_2
XFILLER_0_115_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_204 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17401_ VGND VPWR VPWR VGND _03467_ keymem.key_mem\[14\]\[99\] _03485_ _03486_ sky130_fd_sc_hd__mux2_2
X_11825_ VGND VPWR result[79] _07476_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14613_ VGND VPWR VGND VPWR _10079_ _10077_ _10081_ _10078_ sky130_fd_sc_hd__nand3_2
X_18381_ VPWR VGND VGND VPWR _04274_ _04275_ _04190_ sky130_fd_sc_hd__nor2_2
X_15593_ VGND VPWR VPWR VGND _11051_ keymem.prev_key1_reg\[78\] _11045_ _11046_ _10378_
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_16_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14544_ VPWR VGND VPWR VGND _10007_ _10011_ _10009_ _10005_ _10012_ sky130_fd_sc_hd__or4_2
XFILLER_0_200_377 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17332_ VPWR VGND VGND VPWR keylen _03423_ _03424_ _03425_ sky130_fd_sc_hd__nor3_2
X_11756_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[13\] dec_new_block\[45\]
+ _07442_ sky130_fd_sc_hd__mux2_2
XFILLER_0_95_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_172_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_265_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14475_ VPWR VGND VGND VPWR _09124_ _09944_ _09173_ sky130_fd_sc_hd__nor2_2
X_17263_ VGND VPWR VGND VPWR _03363_ _09637_ _03362_ _02475_ sky130_fd_sc_hd__o21a_2
XFILLER_0_165_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11687_ VGND VPWR result[10] _07407_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_102_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_10_1141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19002_ VGND VPWR _04832_ _04616_ _04831_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_16214_ VGND VPWR VGND VPWR _11386_ _11466_ _02379_ _11400_ sky130_fd_sc_hd__a21oi_2
X_13426_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[126\] _07834_ keymem.key_mem\[10\]\[126\]
+ _07909_ _08903_ sky130_fd_sc_hd__a22o_2
X_17194_ VGND VPWR _02342_ _03299_ _03301_ _03300_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_226_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16145_ VGND VPWR VGND VPWR _11390_ _11348_ _11336_ _11246_ _11599_ sky130_fd_sc_hd__a2bb2o_2
X_13357_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[119\] _07872_ keymem.key_mem\[12\]\[119\]
+ _07620_ _08841_ sky130_fd_sc_hd__a22o_2
XFILLER_0_45_1215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_84_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12308_ VGND VPWR enc_block.round_key\[18\] _07892_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_87_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_114_1_Right_715 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16076_ VPWR VGND VPWR VGND _11528_ _11530_ _11529_ _11220_ _11531_ sky130_fd_sc_hd__or4_2
XFILLER_0_126_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13288_ VPWR VGND VPWR VGND _08778_ keymem.key_mem\[9\]\[112\] _07717_ keymem.key_mem\[8\]\[112\]
+ _07929_ _08779_ sky130_fd_sc_hd__a221o_2
X_15027_ VGND VPWR VGND VPWR _10490_ _10478_ _10462_ _10491_ sky130_fd_sc_hd__a21o_2
XFILLER_0_23_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19904_ VGND VPWR VPWR VGND _05361_ keymem.key_mem\[11\]\[108\] _03543_ _05364_ sky130_fd_sc_hd__mux2_2
X_12239_ VPWR VGND VPWR VGND _07828_ keymem.key_mem\[5\]\[13\] _07595_ keymem.key_mem\[8\]\[13\]
+ _07539_ _07829_ sky130_fd_sc_hd__a221o_2
X_19835_ VGND VPWR _05327_ _03287_ _00703_ _05243_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_209_978 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_194_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_263_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_127_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_237_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19766_ VGND VPWR _00670_ _05291_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_120_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16978_ VPWR VGND VPWR VGND _03106_ key[184] _10322_ sky130_fd_sc_hd__or2_2
XFILLER_0_36_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_195_2_Right_267 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_251_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18717_ VPWR VGND VPWR VGND _04575_ _04550_ _04574_ enc_block.block_w1_reg\[29\]
+ _04328_ _00337_ sky130_fd_sc_hd__a221o_2
XFILLER_0_237_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15929_ VGND VPWR _11385_ _11384_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19697_ VGND VPWR _00637_ _05255_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_155_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18648_ VPWR VGND _04514_ enc_block.block_w1_reg\[30\] enc_block.block_w2_reg\[21\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_188_351 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_204_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_188_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_172_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_91_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_384 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18579_ VPWR VGND _04452_ enc_block.block_w2_reg\[23\] enc_block.block_w3_reg\[14\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_4_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20610_ VGND VPWR VPWR VGND _05736_ _03099_ keymem.key_mem\[8\]\[55\] _05739_ sky130_fd_sc_hd__mux2_2
X_21590_ VGND VPWR VPWR VGND _06259_ _09724_ keymem.key_mem\[4\]\[1\] _06261_ sky130_fd_sc_hd__mux2_2
XFILLER_0_7_822 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_131_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20541_ VGND VPWR _01034_ _05702_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_6_354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23260_ VPWR VGND _07146_ _07145_ enc_block.round_key\[5\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_20472_ VGND VPWR _01002_ _05665_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_54_290 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_162_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22211_ VGND VPWR VPWR VGND _06589_ _02893_ keymem.key_mem\[2\]\[34\] _06593_ sky130_fd_sc_hd__mux2_2
XFILLER_0_166_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23191_ VGND VPWR _02303_ _07083_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_43_997 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_207_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22142_ VGND VPWR _01781_ _06556_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_203_1226 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_61_1050 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22073_ VGND VPWR VPWR VGND _06516_ _05029_ keymem.key_mem\[3\]\[98\] _06519_ sky130_fd_sc_hd__mux2_2
X_21024_ VGND VPWR _01259_ _05960_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_215_915 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25832_ VGND VPWR VPWR VGND clk _02325_ reset_n enc_block.block_w3_reg\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_96_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_242_745 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_184_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1046 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22975_ VGND VPWR VGND VPWR _02218_ _06952_ _06916_ keymem.prev_key1_reg\[41\] sky130_fd_sc_hd__o21a_2
X_25763_ keymem.prev_key1_reg\[79\] clk _02256_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_214_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24714_ VGND VPWR VPWR VGND clk _01207_ reset_n keymem.key_mem\[7\]\[67\] sky130_fd_sc_hd__dfrtp_2
X_21926_ VPWR VGND keymem.key_mem\[3\]\[29\] _06441_ _06439_ VPWR VGND sky130_fd_sc_hd__and2_2
X_25694_ keymem.prev_key1_reg\[10\] clk _02187_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_70_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_384 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_74_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24645_ VGND VPWR VPWR VGND clk _01138_ reset_n keymem.key_mem\[8\]\[126\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_194_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21857_ VPWR VGND _08933_ _06401_ _05241_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_84_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20808_ VPWR VGND keymem.key_mem\[7\]\[18\] _05846_ _05844_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_33_1152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24576_ VGND VPWR VPWR VGND clk _01069_ reset_n keymem.key_mem\[8\]\[57\] sky130_fd_sc_hd__dfrtp_2
X_12590_ VGND VPWR _08150_ _07619_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21788_ VGND VPWR VPWR VGND _06355_ _03459_ keymem.key_mem\[4\]\[95\] _06365_ sky130_fd_sc_hd__mux2_2
XFILLER_0_110_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23527_ VGND VPWR VPWR VGND clk _00028_ reset_n keymem.key_mem\[14\]\[16\] sky130_fd_sc_hd__dfrtp_2
X_20739_ VGND VPWR _01128_ _05806_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_147_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_110_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14260_ VGND VPWR _09730_ _09729_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23458_ VGND VPWR VGND VPWR _07323_ _04064_ _07322_ _07321_ sky130_fd_sc_hd__o21a_2
X_13211_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[104\] _07596_ keymem.key_mem\[8\]\[104\]
+ _07752_ _08710_ sky130_fd_sc_hd__a22o_2
XFILLER_0_208_1137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22409_ VGND VPWR VPWR VGND _06696_ keymem.key_mem\[1\]\[0\] _09537_ _06697_ sky130_fd_sc_hd__mux2_2
X_14191_ VGND VPWR VPWR VGND _09211_ _09662_ _09201_ sky130_fd_sc_hd__and2b_2
XFILLER_0_184_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23389_ VGND VPWR _07262_ enc_block.round_key\[18\] _07261_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_249_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13142_ VPWR VGND VPWR VGND _08647_ keymem.key_mem\[12\]\[97\] _07722_ keymem.key_mem\[8\]\[97\]
+ _08265_ _08648_ sky130_fd_sc_hd__a221o_2
X_25128_ VGND VPWR VPWR VGND clk _01621_ reset_n keymem.key_mem\[4\]\[97\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_81_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17950_ VGND VPWR VPWR VGND _03876_ key[235] keymem.prev_key1_reg\[107\] _03898_
+ sky130_fd_sc_hd__mux2_2
X_13073_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[90\] _08577_ _08585_ _08581_ _08586_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_260_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25059_ VGND VPWR VPWR VGND clk _01552_ reset_n keymem.key_mem\[4\]\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_179 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_104_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16901_ VGND VPWR _00060_ _03036_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12024_ VPWR VGND VPWR VGND _07625_ keymem.key_mem\[11\]\[1\] _07600_ keymem.key_mem\[2\]\[1\]
+ _07546_ _07626_ sky130_fd_sc_hd__a221o_2
XFILLER_0_79_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17881_ VGND VPWR VPWR VGND _03836_ _03850_ keymem.prev_key0_reg\[85\] _03851_ sky130_fd_sc_hd__mux2_2
XFILLER_0_121_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19620_ VGND VPWR VPWR VGND _05205_ _05039_ keymem.key_mem\[12\]\[103\] _05213_ sky130_fd_sc_hd__mux2_2
X_16832_ VGND VPWR _00054_ _02973_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_254_1102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_228_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_195_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19551_ VGND VPWR VPWR VGND _05151_ _04983_ keymem.key_mem\[12\]\[70\] _05177_ sky130_fd_sc_hd__mux2_2
XFILLER_0_73_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16763_ VPWR VGND VGND VPWR _02911_ _11456_ _10088_ sky130_fd_sc_hd__nand2_2
X_13975_ VGND VPWR _09447_ _09300_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_191_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18502_ VGND VPWR _04383_ enc_block.block_w3_reg\[15\] enc_block.block_w2_reg\[23\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15714_ VGND VPWR VGND VPWR enc_block.block_w2_reg\[19\] _09269_ _09021_ _11168_
+ _11170_ _11169_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_87_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_981 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_92_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19482_ VGND VPWR VGND VPWR _05140_ keymem.key_mem_we _02924_ _05135_ _00537_ sky130_fd_sc_hd__a31o_2
X_12926_ VGND VPWR VGND VPWR _07778_ keymem.key_mem\[3\]\[76\] _08450_ _08452_ _08453_
+ _08243_ sky130_fd_sc_hd__a2111o_2
X_16694_ VGND VPWR _02847_ keymem.prev_key0_reg\[127\] _02846_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_18433_ VGND VPWR _04320_ enc_block.block_w1_reg\[24\] enc_block.block_w1_reg\[31\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15645_ VPWR VGND VPWR VGND _11102_ _11101_ sky130_fd_sc_hd__inv_2
X_12857_ VGND VPWR _08391_ _07567_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_180_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_201_664 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11808_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[7\] dec_new_block\[71\]
+ _07468_ sky130_fd_sc_hd__mux2_2
X_18364_ VGND VPWR _04259_ enc_block.block_w3_reg\[3\] enc_block.block_w1_reg\[18\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15576_ VGND VPWR _11035_ keymem.prev_key1_reg\[13\] keymem.prev_key1_reg\[45\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
X_12788_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[62\] _07613_ keymem.key_mem\[14\]\[62\]
+ _07744_ _08329_ sky130_fd_sc_hd__a22o_2
XFILLER_0_145_207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_909 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17315_ VGND VPWR VPWR VGND _03384_ keymem.key_mem\[14\]\[89\] _03409_ _03410_ sky130_fd_sc_hd__mux2_2
X_14527_ VGND VPWR VPWR VGND _09052_ _09101_ _09086_ _09995_ sky130_fd_sc_hd__or3_2
X_11739_ VGND VPWR result[36] _07433_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18295_ VPWR VGND VGND VPWR _04197_ _04194_ _04195_ sky130_fd_sc_hd__nand2_2
XFILLER_0_22_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17246_ VGND VPWR VPWR VGND _03296_ keymem.key_mem\[14\]\[82\] _03347_ _03348_ sky130_fd_sc_hd__mux2_2
X_14458_ VGND VPWR _09927_ _09729_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_189_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_836 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_163_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13409_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[124\] _07613_ keymem.key_mem\[12\]\[124\]
+ _07806_ _08888_ sky130_fd_sc_hd__a22o_2
XFILLER_0_4_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17177_ VGND VPWR VGND VPWR _03281_ key[203] _10908_ _09638_ _03286_ _03285_ sky130_fd_sc_hd__a221oi_2
X_14389_ VGND VPWR VPWR VGND _09859_ _09717_ _09856_ _09858_ _09513_ sky130_fd_sc_hd__o31a_2
XFILLER_0_98_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_625 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16128_ VPWR VGND VGND VPWR _11400_ _11219_ _11280_ _11274_ _11582_ _11581_ sky130_fd_sc_hd__o221a_2
XFILLER_0_267_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_1_Right_716 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16059_ VPWR VGND VGND VPWR _11332_ _11329_ _11514_ _11316_ _11370_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_259_1002 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_209_720 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_202_1270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19818_ VGND VPWR VPWR VGND _05314_ keymem.key_mem\[11\]\[67\] _03217_ _05319_ sky130_fd_sc_hd__mux2_2
XFILLER_0_100_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_138_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19749_ VGND VPWR VPWR VGND _05281_ keymem.key_mem\[11\]\[34\] _02894_ _05283_ sky130_fd_sc_hd__mux2_2
XFILLER_0_78_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22760_ VGND VPWR _06844_ _03287_ _02111_ _06839_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_52_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21711_ VGND VPWR VPWR VGND _06319_ _03129_ keymem.key_mem\[4\]\[58\] _06325_ sky130_fd_sc_hd__mux2_2
XFILLER_0_154_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22691_ VGND VPWR _02070_ _06816_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_250_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24430_ VGND VPWR VPWR VGND clk _00923_ reset_n keymem.key_mem\[9\]\[39\] sky130_fd_sc_hd__dfrtp_2
X_21642_ VGND VPWR VPWR VGND _06286_ _02720_ keymem.key_mem\[4\]\[25\] _06289_ sky130_fd_sc_hd__mux2_2
XFILLER_0_176_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24361_ VGND VPWR VPWR VGND clk _00854_ reset_n keymem.key_mem\[10\]\[98\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_170_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21573_ VGND VPWR VPWR VGND _06242_ _03633_ keymem.key_mem\[5\]\[122\] _06251_ sky130_fd_sc_hd__mux2_2
XFILLER_0_69_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23312_ VPWR VGND VGND VPWR _07192_ _07193_ _04095_ sky130_fd_sc_hd__nor2_2
X_20524_ VGND VPWR VPWR VGND _05692_ _11098_ keymem.key_mem\[8\]\[14\] _05694_ sky130_fd_sc_hd__mux2_2
XFILLER_0_244_1304 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24292_ VGND VPWR VPWR VGND clk _00785_ reset_n keymem.key_mem\[10\]\[29\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_7_685 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_62_569 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_209_1446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23243_ VGND VPWR _07130_ enc_block.block_w3_reg\[27\] _07129_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_209_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20455_ VGND VPWR _00994_ _05656_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_43_794 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_127_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23174_ VGND VPWR VPWR VGND _07054_ _07072_ keymem.prev_key1_reg\[120\] _07073_ sky130_fd_sc_hd__mux2_2
X_20386_ VGND VPWR _00961_ _05620_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_179_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22125_ VGND VPWR VPWR VGND _06538_ _05081_ keymem.key_mem\[3\]\[123\] _06546_ sky130_fd_sc_hd__mux2_2
XFILLER_0_30_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_321 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_247_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_112_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_499 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22056_ VPWR VGND keymem.key_mem\[3\]\[90\] _06510_ _06484_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_220_1381 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21007_ VGND VPWR _01251_ _05951_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_199_402 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25815_ VGND VPWR VPWR VGND clk _02308_ reset_n enc_block.block_w3_reg\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_230_704 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_230_715 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_138_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13760_ VGND VPWR VGND VPWR _09053_ _09056_ _09077_ _09040_ _09071_ _09232_ sky130_fd_sc_hd__o32a_2
X_22958_ VGND VPWR VGND VPWR _02898_ _03794_ _02902_ _06942_ sky130_fd_sc_hd__a21o_2
X_25746_ keymem.prev_key1_reg\[62\] clk _02239_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_69_146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_74_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_165_1_Left_432 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12711_ VGND VPWR _08259_ _07534_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21909_ VGND VPWR VGND VPWR _06431_ keymem.key_mem_we _02550_ _06420_ _01673_ sky130_fd_sc_hd__a31o_2
X_13691_ VGND VPWR VGND VPWR _09163_ _09162_ _09161_ _09158_ _09155_ sky130_fd_sc_hd__and4_2
XFILLER_0_84_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25677_ VGND VPWR VPWR VGND clk _02170_ reset_n keymem.rcon_logic.tmp_rcon\[7\] sky130_fd_sc_hd__dfrtp_2
X_22889_ VGND VPWR _02185_ _06899_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_84_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_133_2_Left_604 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15430_ VPWR VGND VPWR VGND _10889_ _10890_ _10891_ _10882_ _10884_ sky130_fd_sc_hd__or4b_2
X_12642_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[48\] _07579_ keymem.key_mem\[8\]\[48\]
+ _07878_ _08197_ sky130_fd_sc_hd__a22o_2
XFILLER_0_38_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24628_ VGND VPWR VPWR VGND clk _01121_ reset_n keymem.key_mem\[8\]\[109\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_127_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_182_302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15361_ VPWR VGND VPWR VGND _10823_ keymem.prev_key0_reg\[10\] sky130_fd_sc_hd__inv_2
X_12573_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[41\] _08124_ _08134_ _08129_ enc_block.round_key\[41\]
+ sky130_fd_sc_hd__o22a_2
X_24559_ VGND VPWR VPWR VGND clk _01052_ reset_n keymem.key_mem\[8\]\[40\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_1201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17100_ VGND VPWR _03217_ _03216_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14312_ VGND VPWR VGND VPWR _09327_ _09582_ _09749_ _09375_ _09782_ sky130_fd_sc_hd__o22a_2
XPHY_EDGE_ROW_158_2_Right_230 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15292_ VGND VPWR VGND VPWR _10569_ _10538_ _10754_ _10668_ sky130_fd_sc_hd__a21oi_2
X_18080_ VPWR VGND VPWR VGND _04000_ _03996_ _03998_ sky130_fd_sc_hd__or2_2
XFILLER_0_227_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_262 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14243_ VPWR VGND VPWR VGND _09712_ _09714_ _09710_ _09711_ sky130_fd_sc_hd__or3b_2
X_17031_ VPWR VGND VPWR VGND _03154_ key[61] _09719_ sky130_fd_sc_hd__or2_2
XFILLER_0_0_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_145_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14174_ VGND VPWR VPWR VGND _09108_ _09082_ _09189_ _09645_ sky130_fd_sc_hd__or3_2
XFILLER_0_106_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_145_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13125_ VGND VPWR enc_block.round_key\[95\] _08632_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18982_ VPWR VGND VPWR VGND _04814_ _04788_ _04813_ enc_block.block_w2_reg\[23\]
+ _04709_ _00363_ sky130_fd_sc_hd__a221o_2
X_17933_ VGND VPWR _00242_ _03886_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13056_ VPWR VGND VPWR VGND _08569_ keymem.key_mem\[11\]\[89\] _07781_ keymem.key_mem\[2\]\[89\]
+ _07698_ _08570_ sky130_fd_sc_hd__a221o_2
XFILLER_0_264_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_206_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12007_ VGND VPWR _07609_ _07608_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_246_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17864_ VGND VPWR _00220_ _03839_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_128_2_Left_599 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19603_ VPWR VGND keymem.key_mem\[12\]\[95\] _05204_ _05094_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_255_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16815_ VGND VPWR VGND VPWR _02957_ _02342_ _02958_ _10664_ sky130_fd_sc_hd__nand3_2
XFILLER_0_156_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_219_1052 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17795_ VGND VPWR _03792_ _10371_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_191_1244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_97_1_Left_364 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19534_ VPWR VGND keymem.key_mem\[12\]\[62\] _05168_ _05158_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_156_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16746_ VGND VPWR _00046_ _02895_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13958_ VPWR VGND VPWR VGND _09307_ _09309_ _09339_ _09338_ _09430_ sky130_fd_sc_hd__or4_2
XFILLER_0_92_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_2_Left_536 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_117_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19465_ VPWR VGND keymem.key_mem\[12\]\[30\] _05131_ _05128_ VPWR VGND sky130_fd_sc_hd__and2_2
X_12909_ VGND VPWR VGND VPWR _08438_ _07712_ keymem.key_mem\[6\]\[74\] _08435_ _08437_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_5_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16677_ VGND VPWR VGND VPWR _02829_ _02828_ _02830_ _02831_ sky130_fd_sc_hd__a21o_2
XFILLER_0_9_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13889_ VGND VPWR _09361_ _09315_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_53_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18416_ enc_block.sword_ctr_reg\[1\] _04305_ _08945_ _03972_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__and3_2
XFILLER_0_75_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_235_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_472 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_140 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15628_ VGND VPWR VGND VPWR _10513_ _10522_ _10867_ _10633_ _10580_ _11086_ sky130_fd_sc_hd__o32a_2
XFILLER_0_8_405 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1304 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19396_ VGND VPWR _05092_ _05091_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18347_ VPWR VGND VPWR VGND _04244_ _04162_ _04242_ sky130_fd_sc_hd__or2_2
XFILLER_0_5_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15559_ VPWR VGND VPWR VGND _11005_ _11017_ _11010_ _10995_ _11018_ sky130_fd_sc_hd__or4_2
XFILLER_0_44_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_189_1195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_558 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18278_ VPWR VGND _04181_ enc_block.block_w2_reg\[10\] enc_block.block_w3_reg\[3\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_140_43 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_86_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17229_ VPWR VGND VPWR VGND _03332_ keymem.prev_key0_reg\[81\] sky130_fd_sc_hd__inv_2
XFILLER_0_163_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_934 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_25_794 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20240_ VGND VPWR VPWR VGND _05535_ _10662_ keymem.key_mem\[9\]\[8\] _05544_ sky130_fd_sc_hd__mux2_2
XFILLER_0_124_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_163_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20171_ VGND VPWR VPWR VGND _05504_ _03525_ keymem.key_mem\[10\]\[105\] _05506_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_116_1_Right_717 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_120_2_Right_192 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_196_1111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_149_96 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23930_ VGND VPWR VPWR VGND clk _00423_ reset_n keymem.key_mem\[13\]\[51\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1130 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23861_ VGND VPWR VPWR VGND clk _00354_ reset_n enc_block.block_w2_reg\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_174_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25600_ VGND VPWR VPWR VGND clk _02093_ reset_n keymem.key_mem\[0\]\[57\] sky130_fd_sc_hd__dfrtp_2
X_22812_ VGND VPWR _06860_ _06779_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_174_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23792_ VGND VPWR VPWR VGND clk _00285_ reset_n enc_block.block_w0_reg\[11\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_71_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_75_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_135_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22743_ VGND VPWR _06837_ _06779_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25531_ VGND VPWR VPWR VGND clk _02024_ reset_n keymem.key_mem\[1\]\[116\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_71_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25462_ VGND VPWR VPWR VGND clk _01955_ reset_n keymem.key_mem\[1\]\[47\] sky130_fd_sc_hd__dfrtp_2
X_22674_ VGND VPWR _02061_ _06808_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_164_302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24413_ VGND VPWR VPWR VGND clk _00906_ reset_n keymem.key_mem\[9\]\[22\] sky130_fd_sc_hd__dfrtp_2
X_21625_ VGND VPWR VPWR VGND _06275_ _11546_ keymem.key_mem\[4\]\[17\] _06280_ sky130_fd_sc_hd__mux2_2
X_25393_ VGND VPWR VPWR VGND clk _01886_ reset_n keymem.key_mem\[2\]\[106\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_8_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24344_ VGND VPWR VPWR VGND clk _00837_ reset_n keymem.key_mem\[10\]\[81\] sky130_fd_sc_hd__dfrtp_2
X_21556_ VGND VPWR _06242_ _06115_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_63_867 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20507_ VGND VPWR VPWR VGND _05680_ _10283_ keymem.key_mem\[8\]\[6\] _05685_ sky130_fd_sc_hd__mux2_2
XFILLER_0_181_1413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_62_377 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24275_ VGND VPWR VPWR VGND clk _00768_ reset_n keymem.key_mem\[10\]\[12\] sky130_fd_sc_hd__dfrtp_2
X_21487_ VGND VPWR VPWR VGND _06196_ _03339_ keymem.key_mem\[5\]\[81\] _06206_ sky130_fd_sc_hd__mux2_2
XFILLER_0_181_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23226_ VGND VPWR _07114_ _04005_ _02307_ _07096_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_82_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20438_ VGND VPWR _00986_ _05647_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_142_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_753 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_43_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_181_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_775 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_261_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23157_ VGND VPWR VPWR VGND _07054_ _03572_ keymem.prev_key1_reg\[113\] _07063_ sky130_fd_sc_hd__mux2_2
XFILLER_0_31_797 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_43_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20369_ VGND VPWR _00953_ _05611_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_222_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22108_ VGND VPWR VPWR VGND _06527_ _05064_ keymem.key_mem\[3\]\[115\] _06537_ sky130_fd_sc_hd__mux2_2
XFILLER_0_100_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23088_ VGND VPWR VPWR VGND _02264_ _03387_ _03391_ _06976_ _07019_ sky130_fd_sc_hd__o31a_2
X_14930_ VGND VPWR VGND VPWR _10394_ enc_block.block_w2_reg\[8\] enc_block.sword_ctr_reg\[1\]
+ enc_block.sword_ctr_reg\[0\] sky130_fd_sc_hd__and3b_2
X_22039_ VGND VPWR _01733_ _06501_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_261_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14861_ key[135] _10326_ keylen _10325_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_243_873 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16600_ VGND VPWR VGND VPWR _02756_ _02755_ keymem.prev_key1_reg\[91\] _02757_ sky130_fd_sc_hd__a21o_2
X_13812_ VPWR VGND VPWR VGND _09284_ enc_block.block_w0_reg\[29\] _08952_ sky130_fd_sc_hd__or2_2
XFILLER_0_153_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17580_ VGND VPWR VPWR VGND _03593_ keymem.key_mem\[14\]\[123\] _03640_ _03641_ sky130_fd_sc_hd__mux2_2
XFILLER_0_192_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14792_ VGND VPWR VGND VPWR _09563_ _09352_ _09559_ _10258_ sky130_fd_sc_hd__a21o_2
XFILLER_0_216_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_1000 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16531_ VGND VPWR _00036_ _02690_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_153_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13743_ VPWR VGND VPWR VGND _09215_ _09089_ sky130_fd_sc_hd__inv_2
X_25729_ keymem.prev_key1_reg\[45\] clk _02222_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_35_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_230_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19250_ VGND VPWR _00449_ _04996_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_211_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16462_ VGND VPWR VGND VPWR _11336_ _11282_ _11252_ _11385_ _02623_ sky130_fd_sc_hd__o22a_2
XFILLER_0_70_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13674_ VGND VPWR _09146_ _09145_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_6_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18201_ VGND VPWR _04111_ _04022_ _04110_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_210_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_110 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15413_ VPWR VGND VPWR VGND _10865_ _10873_ _10869_ _10676_ _10874_ sky130_fd_sc_hd__or4_2
XFILLER_0_2_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12625_ VGND VPWR VGND VPWR _07536_ keymem.key_mem\[0\]\[46\] _08181_ _08176_ _08174_
+ _08182_ sky130_fd_sc_hd__o32a_2
X_19181_ VPWR VGND keymem.key_mem_we _04955_ _03056_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16393_ VGND VPWR VGND VPWR _02555_ _11311_ _11380_ _11306_ _11460_ _11239_ sky130_fd_sc_hd__a41o_2
X_18132_ VPWR VGND VPWR VGND _04048_ _04044_ _04046_ sky130_fd_sc_hd__or2_2
X_15344_ VPWR VGND VPWR VGND _10803_ _10805_ _10804_ _10802_ _10806_ sky130_fd_sc_hd__or4_2
X_12556_ VGND VPWR VGND VPWR _07731_ keymem.key_mem\[13\]\[40\] _08115_ _08118_ _08119_
+ _07574_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_53_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_80_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_159_2_Right_231 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18063_ VGND VPWR _03984_ enc_block.block_w2_reg\[9\] _03960_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_12487_ VGND VPWR enc_block.round_key\[33\] _08056_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15275_ _09679_ _10738_ keymem.prev_key1_reg\[105\] _09708_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_17014_ VPWR VGND VPWR VGND _03138_ _02677_ _03133_ key[187] _02723_ _03139_ sky130_fd_sc_hd__a221o_2
X_14226_ VPWR VGND VGND VPWR _09696_ _09697_ _09692_ sky130_fd_sc_hd__nor2_2
XFILLER_0_262_1278 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_223_1229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_160_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14157_ VPWR VGND VPWR VGND _09615_ _09627_ _09620_ _09610_ _09628_ sky130_fd_sc_hd__or4_2
XFILLER_0_201_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_240_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_119_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13108_ VPWR VGND VPWR VGND _08616_ keymem.key_mem\[5\]\[94\] _07811_ keymem.key_mem\[13\]\[94\]
+ _07622_ _08617_ sky130_fd_sc_hd__a221o_2
X_14088_ VGND VPWR _09559_ _09335_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18965_ VPWR VGND _04799_ enc_block.block_w0_reg\[13\] enc_block.block_w1_reg\[6\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_201_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17916_ VGND VPWR VPWR VGND _03874_ _03873_ keymem.prev_key0_reg\[96\] _03875_ sky130_fd_sc_hd__mux2_2
X_13039_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[87\] _07674_ keymem.key_mem\[1\]\[87\]
+ _07670_ _08555_ sky130_fd_sc_hd__a22o_2
XFILLER_0_185_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18896_ VGND VPWR _04737_ enc_block.block_w1_reg\[6\] enc_block.block_w1_reg\[7\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17847_ VGND VPWR VPWR VGND _03814_ _03827_ keymem.prev_key0_reg\[74\] _03828_ sky130_fd_sc_hd__mux2_2
XFILLER_0_135_21 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17778_ VGND VPWR _00193_ _03780_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_44_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1145 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_221_545 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19517_ VPWR VGND keymem.key_mem\[12\]\[54\] _05159_ _05158_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_49_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16729_ VGND VPWR VPWR VGND _09511_ key[161] keymem.prev_key1_reg\[33\] _02880_ sky130_fd_sc_hd__mux2_2
XFILLER_0_92_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19448_ VPWR VGND keymem.key_mem\[12\]\[22\] _05122_ _05116_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_18_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_352 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_88_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_363 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19379_ VGND VPWR _00494_ _05080_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21410_ VGND VPWR VPWR VGND _06162_ _02998_ keymem.key_mem\[5\]\[44\] _06166_ sky130_fd_sc_hd__mux2_2
XFILLER_0_151_75 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_263_1009 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22390_ VGND VPWR _01899_ _06686_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_44_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21341_ VPWR VGND VGND VPWR _06130_ keymem.key_mem\[5\]\[11\] _06114_ sky130_fd_sc_hd__nand2_2
XFILLER_0_71_174 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_4_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24060_ VGND VPWR VPWR VGND clk _00553_ reset_n keymem.key_mem\[12\]\[53\] sky130_fd_sc_hd__dfrtp_2
X_21272_ VGND VPWR VPWR VGND _06087_ _03543_ keymem.key_mem\[6\]\[108\] _06092_ sky130_fd_sc_hd__mux2_2
XFILLER_0_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23011_ VPWR VGND VPWR VGND _06974_ keymem.prev_key1_reg\[56\] _06926_ sky130_fd_sc_hd__or2_2
XFILLER_0_64_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20223_ VGND VPWR _05535_ _05534_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_29_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_69_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1217 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_60_1126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20154_ VGND VPWR VPWR VGND _05493_ _03474_ keymem.key_mem\[10\]\[97\] _05497_ sky130_fd_sc_hd__mux2_2
XFILLER_0_244_604 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_99_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_1_Right_718 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_121_2_Right_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24962_ VGND VPWR VPWR VGND clk _01455_ reset_n keymem.key_mem\[5\]\[59\] sky130_fd_sc_hd__dfrtp_2
X_20085_ VGND VPWR VPWR VGND _05457_ _03194_ keymem.key_mem\[10\]\[64\] _05461_ sky130_fd_sc_hd__mux2_2
XFILLER_0_176_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23913_ VGND VPWR VPWR VGND clk _00406_ reset_n keymem.key_mem\[13\]\[34\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24893_ VGND VPWR VPWR VGND clk _01386_ reset_n keymem.key_mem\[6\]\[118\] sky130_fd_sc_hd__dfrtp_2
X_23844_ VGND VPWR VPWR VGND clk _00337_ reset_n enc_block.block_w1_reg\[29\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_135_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_252 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_254_Right_123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23775_ VGND VPWR VPWR VGND clk _00001_ reset_n enc_block.enc_ctrl_reg\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_75_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20987_ VGND VPWR VPWR VGND _05934_ _05037_ keymem.key_mem\[7\]\[102\] _05941_ sky130_fd_sc_hd__mux2_2
XFILLER_0_71_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25514_ VGND VPWR VPWR VGND clk _02007_ reset_n keymem.key_mem\[1\]\[99\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_233 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22726_ VGND VPWR VPWR VGND _06822_ keymem.key_mem\[0\]\[58\] _03130_ _06828_ sky130_fd_sc_hd__mux2_2
XFILLER_0_36_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_211_1133 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_54_108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25445_ VGND VPWR VPWR VGND clk _01938_ reset_n keymem.key_mem\[1\]\[30\] sky130_fd_sc_hd__dfrtp_2
X_22657_ VGND VPWR VPWR VGND _06798_ keymem.key_mem\[0\]\[17\] _11547_ _06800_ sky130_fd_sc_hd__mux2_2
XFILLER_0_211_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12410_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[27\] _07577_ keymem.key_mem\[4\]\[27\]
+ _07550_ _07986_ sky130_fd_sc_hd__a22o_2
X_21608_ VGND VPWR VPWR VGND _06263_ _10746_ keymem.key_mem\[4\]\[9\] _06271_ sky130_fd_sc_hd__mux2_2
X_13390_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[122\] _08216_ keymem.key_mem\[8\]\[122\]
+ _07541_ _08871_ sky130_fd_sc_hd__a22o_2
XFILLER_0_63_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25376_ VGND VPWR VPWR VGND clk _01869_ reset_n keymem.key_mem\[2\]\[89\] sky130_fd_sc_hd__dfrtp_2
X_22588_ VGND VPWR _06774_ _03859_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12341_ VGND VPWR enc_block.round_key\[20\] _07923_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24327_ VGND VPWR VPWR VGND clk _00820_ reset_n keymem.key_mem\[10\]\[64\] sky130_fd_sc_hd__dfrtp_2
X_21539_ VGND VPWR _01501_ _06233_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_51_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_580 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_107_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15060_ VPWR VGND VPWR VGND _10483_ _10477_ _10440_ _10451_ _10524_ sky130_fd_sc_hd__or4_2
X_24258_ VGND VPWR VPWR VGND clk _00751_ reset_n keymem.key_mem\[11\]\[123\] sky130_fd_sc_hd__dfrtp_2
X_12272_ VGND VPWR enc_block.round_key\[15\] _07859_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_146_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14011_ VGND VPWR VGND VPWR _09473_ _09472_ _09477_ _09481_ _09483_ _09482_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_82_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23209_ VPWR VGND _07099_ enc_block.block_w0_reg\[17\] enc_block.block_w3_reg\[25\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_47_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24189_ VGND VPWR VPWR VGND clk _00682_ reset_n keymem.key_mem\[11\]\[54\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_82_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1251 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_219_122 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_43_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18750_ VGND VPWR _04605_ enc_block.block_w2_reg\[24\] _04604_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15962_ _11340_ _11418_ _11258_ _11417_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_179_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17701_ VGND VPWR _03732_ _02647_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14913_ VPWR VGND _10375_ _10377_ _10376_ VPWR VGND sky130_fd_sc_hd__and2_2
X_18681_ VGND VPWR _04543_ _03977_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_222_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15893_ VGND VPWR VGND VPWR _11349_ _11221_ _11286_ _11174_ _11263_ sky130_fd_sc_hd__and4_2
XFILLER_0_236_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_810 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17632_ VGND VPWR VPWR VGND _03681_ _03683_ keymem.prev_key0_reg\[3\] _03684_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_262_Left_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14844_ VGND VPWR VGND VPWR _09343_ _09411_ _09397_ _09419_ _10309_ sky130_fd_sc_hd__o22a_2
XFILLER_0_153_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_114_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17563_ VPWR VGND VGND VPWR keylen _03624_ _03625_ _03626_ sky130_fd_sc_hd__nor3_2
X_14775_ VPWR VGND VGND VPWR _09450_ _09350_ _09381_ _09386_ _10241_ _10240_ sky130_fd_sc_hd__o221a_2
XFILLER_0_93_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_948 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_85_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11987_ VPWR VGND VGND VPWR _07537_ _07590_ _07554_ sky130_fd_sc_hd__nor2_2
X_19302_ VGND VPWR _00469_ _05028_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_252_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16514_ VGND VPWR _02674_ keymem.prev_key0_reg\[24\] _02673_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_13726_ VPWR VGND VGND VPWR _09195_ _09197_ _09198_ sky130_fd_sc_hd__or2b_2
XFILLER_0_15_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_188_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17494_ VPWR VGND VGND VPWR _03565_ _03566_ keylen sky130_fd_sc_hd__nor2_2
XFILLER_0_54_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19233_ VGND VPWR VGND VPWR _04985_ keymem.key_mem_we _03252_ _04968_ _00443_ sky130_fd_sc_hd__a31o_2
XFILLER_0_252_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16445_ VPWR VGND VPWR VGND _02606_ _10085_ _02596_ key[150] _11043_ _02607_ sky130_fd_sc_hd__a221o_2
X_13657_ VGND VPWR VPWR VGND _09058_ _09039_ _09057_ _09129_ sky130_fd_sc_hd__or3_2
XFILLER_0_128_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_264_1307 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19164_ VGND VPWR VPWR VGND _04928_ _04943_ keymem.key_mem\[13\]\[44\] _04944_ sky130_fd_sc_hd__mux2_2
X_12608_ VPWR VGND VPWR VGND _08165_ keymem.key_mem\[10\]\[45\] _07562_ keymem.key_mem\[12\]\[45\]
+ _07894_ _08166_ sky130_fd_sc_hd__a221o_2
X_16376_ VGND VPWR VGND VPWR _02539_ _02538_ _02537_ keymem.prev_key0_reg\[117\] sky130_fd_sc_hd__and3b_2
X_13588_ VPWR VGND VGND VPWR _09060_ _09051_ _09039_ sky130_fd_sc_hd__nand2_2
XFILLER_0_264_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_143_327 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_121_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18115_ VGND VPWR _04032_ enc_block.block_w2_reg\[13\] enc_block.block_w1_reg\[21\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15327_ VPWR VGND VPWR VGND _10787_ _10788_ _10789_ _10701_ _10786_ sky130_fd_sc_hd__or4b_2
XFILLER_0_42_826 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_54_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12539_ VGND VPWR VGND VPWR _07737_ keymem.key_mem\[1\]\[38\] _08100_ _08102_ _08104_
+ _08103_ sky130_fd_sc_hd__a2111o_2
X_19095_ VPWR VGND keymem.key_mem\[13\]\[17\] _04902_ _04887_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_30_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18046_ VPWR VGND VPWR VGND _03967_ block[96] _03959_ enc_block.block_w3_reg\[0\]
+ _03954_ _03968_ sky130_fd_sc_hd__a221o_2
XFILLER_0_227_1173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15258_ VPWR VGND VGND VPWR _10611_ _10721_ _10573_ sky130_fd_sc_hd__nor2_2
XFILLER_0_129_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_164_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1_444 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14209_ VGND VPWR VGND VPWR _09210_ _09145_ _09016_ _09072_ _09680_ sky130_fd_sc_hd__o22a_2
XFILLER_0_61_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15189_ VPWR VGND _10552_ _10653_ _10652_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_199_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_61_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_205_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19997_ VGND VPWR VPWR VGND _05413_ _02608_ keymem.key_mem\[10\]\[22\] _05415_ sky130_fd_sc_hd__mux2_2
XFILLER_0_123_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_254_946 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18948_ VGND VPWR _04784_ _04781_ _04783_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_18879_ VGND VPWR VGND VPWR _04720_ _04719_ _04722_ _04718_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_101_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20910_ VGND VPWR VPWR VGND _05880_ _04975_ keymem.key_mem\[7\]\[65\] _05901_ sky130_fd_sc_hd__mux2_2
XFILLER_0_262_990 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_238_1280 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21890_ VGND VPWR VGND VPWR _06421_ keymem.key_mem_we _10977_ _06420_ _01664_ sky130_fd_sc_hd__a31o_2
XFILLER_0_171_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20841_ VGND VPWR _01173_ _05863_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_72_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23560_ VGND VPWR VPWR VGND clk _00061_ reset_n keymem.key_mem\[14\]\[49\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20772_ VGND VPWR VGND VPWR _05826_ keymem.key_mem_we _09725_ _05821_ _01141_ sky130_fd_sc_hd__a31o_2
XFILLER_0_33_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_266 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22511_ VGND VPWR VPWR VGND _06739_ keymem.key_mem\[1\]\[56\] _03109_ _06743_ sky130_fd_sc_hd__mux2_2
X_23491_ VGND VPWR _07352_ _07149_ _07351_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_247_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_212_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_112_1_Left_379 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25230_ VGND VPWR VPWR VGND clk _01723_ reset_n keymem.key_mem\[3\]\[71\] sky130_fd_sc_hd__dfrtp_2
X_22442_ VGND VPWR _01923_ _06714_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_146_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_601 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_826 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25161_ VGND VPWR VPWR VGND clk _01654_ reset_n keymem.key_mem\[3\]\[2\] sky130_fd_sc_hd__dfrtp_2
X_22373_ VGND VPWR _01891_ _06677_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_32_336 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_60_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24112_ VGND VPWR VPWR VGND clk _00605_ reset_n keymem.key_mem\[12\]\[105\] sky130_fd_sc_hd__dfrtp_2
X_21324_ VGND VPWR VPWR VGND _06117_ _09991_ keymem.key_mem\[5\]\[3\] _06121_ sky130_fd_sc_hd__mux2_2
XFILLER_0_143_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25092_ VGND VPWR VPWR VGND clk _01585_ reset_n keymem.key_mem\[4\]\[61\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_182_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1284 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24043_ VGND VPWR VPWR VGND clk _00536_ reset_n keymem.key_mem\[12\]\[36\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_143_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21255_ VGND VPWR VPWR VGND _06076_ _03492_ keymem.key_mem\[6\]\[100\] _06083_ sky130_fd_sc_hd__mux2_2
XFILLER_0_241_1159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_198_1003 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_229_431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_174_1_Left_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20206_ VGND VPWR VPWR VGND _05515_ _03633_ keymem.key_mem\[10\]\[122\] _05524_ sky130_fd_sc_hd__mux2_2
X_21186_ VGND VPWR VPWR VGND _06040_ _03216_ keymem.key_mem\[6\]\[67\] _06047_ sky130_fd_sc_hd__mux2_2
XFILLER_0_245_913 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_142_2_Left_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_245_946 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20137_ VGND VPWR VPWR VGND _05482_ _03409_ keymem.key_mem\[10\]\[89\] _05488_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_118_1_Right_719 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_122_2_Right_194 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_254_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20068_ VGND VPWR VPWR VGND _05446_ _03109_ keymem.key_mem\[10\]\[56\] _05452_ sky130_fd_sc_hd__mux2_2
X_24945_ VGND VPWR VPWR VGND clk _01438_ reset_n keymem.key_mem\[5\]\[42\] sky130_fd_sc_hd__dfrtp_2
X_11910_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[26\] dec_new_block\[122\]
+ _07519_ sky130_fd_sc_hd__mux2_2
X_24876_ VGND VPWR VPWR VGND clk _01369_ reset_n keymem.key_mem\[6\]\[101\] sky130_fd_sc_hd__dfrtp_2
X_12890_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[72\] _08124_ _08420_ _08416_ _08421_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_212_320 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_213_1206 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11841_ VGND VPWR result[87] _07484_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23827_ VGND VPWR VPWR VGND clk _00320_ reset_n enc_block.block_w1_reg\[12\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_150_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_200_526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14560_ VGND VPWR VGND VPWR _09146_ _09125_ _09128_ _09140_ _10028_ sky130_fd_sc_hd__o22a_2
X_11772_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[21\] dec_new_block\[53\]
+ _07450_ sky130_fd_sc_hd__mux2_2
X_23758_ keymem.prev_key0_reg\[114\] clk _00255_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_230_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13511_ VGND VPWR _08983_ _08941_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_67_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22709_ VGND VPWR _02083_ _06821_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14491_ VPWR VGND VPWR VGND _09958_ _09959_ _09960_ _09218_ _09957_ sky130_fd_sc_hd__or4b_2
X_23689_ keymem.prev_key0_reg\[45\] clk _00186_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_3_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16230_ VGND VPWR VPWR VGND keymem.round_ctr_reg\[0\] _02394_ _02344_ _02395_ sky130_fd_sc_hd__mux2_2
X_13442_ VPWR VGND VPWR VGND _08917_ keymem.key_mem\[13\]\[127\] _08125_ keymem.key_mem\[12\]\[127\]
+ _07894_ _08918_ sky130_fd_sc_hd__a221o_2
X_25428_ VGND VPWR VPWR VGND clk _01921_ reset_n keymem.key_mem\[1\]\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_137_187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_709 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16161_ VPWR VGND VPWR VGND _11613_ _11614_ _11615_ _11611_ _11612_ sky130_fd_sc_hd__or4b_2
X_13373_ VGND VPWR VGND VPWR _08856_ _07731_ keymem.key_mem\[13\]\[120\] _08853_ _08855_
+ sky130_fd_sc_hd__a211o_2
X_25359_ VGND VPWR VPWR VGND clk _01852_ reset_n keymem.key_mem\[2\]\[72\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_859 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15112_ VGND VPWR VGND VPWR _10543_ _10536_ _10575_ _10574_ _10576_ sky130_fd_sc_hd__o22a_2
X_12324_ VGND VPWR enc_block.round_key\[19\] _07907_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16092_ VGND VPWR _11547_ _11546_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_133_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15043_ VGND VPWR _10507_ _10506_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12255_ VGND VPWR _07844_ _07843_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19920_ VGND VPWR _05372_ _05242_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_74_2_Left_545 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19851_ VGND VPWR VPWR VGND _05328_ keymem.key_mem\[11\]\[83\] _03356_ _05336_ sky130_fd_sc_hd__mux2_2
XFILLER_0_107_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12186_ VGND VPWR _07779_ _07613_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18802_ VPWR VGND _04653_ _04652_ enc_block.round_key\[37\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_208_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_257_1111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19782_ VGND VPWR VPWR VGND _05292_ keymem.key_mem\[11\]\[50\] _03056_ _05300_ sky130_fd_sc_hd__mux2_2
X_16994_ VGND VPWR _00069_ _03120_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_78_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18733_ VPWR VGND VGND VPWR _04316_ _04590_ _04301_ sky130_fd_sc_hd__nor2_2
XFILLER_0_247_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15945_ VGND VPWR VGND VPWR _11397_ _11296_ _11401_ _11400_ sky130_fd_sc_hd__a21oi_2
X_18664_ VPWR VGND VPWR VGND _04528_ _04459_ _04527_ enc_block.block_w1_reg\[23\]
+ _04424_ _00331_ sky130_fd_sc_hd__a221o_2
XFILLER_0_262_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15876_ VGND VPWR _11332_ _11331_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17615_ VGND VPWR _03670_ _10371_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_118_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14827_ VGND VPWR VGND VPWR _10060_ _10292_ _10247_ _10291_ _10107_ sky130_fd_sc_hd__and4bb_2
X_18595_ VGND VPWR _04467_ enc_block.round_key\[80\] _04466_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_231_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_59_734 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_391 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_118_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17546_ VGND VPWR VPWR VGND _10378_ _03610_ key[247] _03611_ sky130_fd_sc_hd__mux2_2
XFILLER_0_148_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14758_ VGND VPWR VGND VPWR _09083_ _09160_ _10224_ _09178_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_58_244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_59_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_929 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_15_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13709_ VGND VPWR _09181_ _09086_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17477_ VGND VPWR _00121_ _03551_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14689_ VPWR VGND VPWR VGND _10148_ _10155_ _10151_ _09206_ _10156_ sky130_fd_sc_hd__or4_2
XFILLER_0_73_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19216_ VPWR VGND keymem.key_mem_we _04975_ _03202_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16428_ VGND VPWR _02590_ keymem.prev_key0_reg\[54\] keymem.prev_key0_reg\[86\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_327 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19147_ VGND VPWR _00410_ _04932_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16359_ VGND VPWR VGND VPWR _11246_ _11204_ _11182_ _11370_ _02522_ sky130_fd_sc_hd__o22a_2
XFILLER_0_15_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_124_360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19078_ VGND VPWR VGND VPWR _04892_ keymem.key_mem_we _10747_ _04878_ _00381_ sky130_fd_sc_hd__a31o_2
XFILLER_0_125_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18029_ VGND VPWR _03951_ _03950_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_41_188 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_125_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21040_ VGND VPWR _01267_ _05968_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_22_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_564 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_732 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_199_1389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_96_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1091 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22991_ VGND VPWR VGND VPWR _02224_ _06962_ _06954_ keymem.prev_key1_reg\[47\] sky130_fd_sc_hd__o21a_2
XFILLER_0_226_489 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24730_ VGND VPWR VPWR VGND clk _01223_ reset_n keymem.key_mem\[7\]\[83\] sky130_fd_sc_hd__dfrtp_2
X_21942_ VGND VPWR VPWR VGND _06449_ _04927_ keymem.key_mem\[3\]\[36\] _06450_ sky130_fd_sc_hd__mux2_2
XFILLER_0_206_180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_136_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24661_ VGND VPWR VPWR VGND clk _01154_ reset_n keymem.key_mem\[7\]\[14\] sky130_fd_sc_hd__dfrtp_2
X_21873_ VPWR VGND keymem.key_mem\[3\]\[5\] _06412_ _06406_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_166_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23612_ VGND VPWR VPWR VGND clk _00113_ reset_n keymem.key_mem\[14\]\[101\] sky130_fd_sc_hd__dfrtp_2
X_20824_ VGND VPWR VGND VPWR _05854_ keymem.key_mem_we _02721_ _05850_ _01165_ sky130_fd_sc_hd__a31o_2
XFILLER_0_136_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24592_ VGND VPWR VPWR VGND clk _01085_ reset_n keymem.key_mem\[8\]\[73\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20755_ VGND VPWR _01136_ _05814_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23543_ VGND VPWR VPWR VGND clk _00044_ reset_n keymem.key_mem\[14\]\[32\] sky130_fd_sc_hd__dfrtp_2
X_23474_ VPWR VGND VGND VPWR _07337_ _07130_ _07336_ sky130_fd_sc_hd__nand2_2
XFILLER_0_68_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20686_ VGND VPWR _01103_ _05778_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25213_ VGND VPWR VPWR VGND clk _01706_ reset_n keymem.key_mem\[3\]\[54\] sky130_fd_sc_hd__dfrtp_2
X_22425_ VGND VPWR _06706_ _03859_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_208_1308 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22356_ VGND VPWR _01883_ _06668_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25144_ VGND VPWR VPWR VGND clk _01637_ reset_n keymem.key_mem\[4\]\[113\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_108_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_147_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21307_ VGND VPWR VPWR VGND _05971_ _03654_ keymem.key_mem\[6\]\[125\] _06110_ sky130_fd_sc_hd__mux2_2
X_25075_ VGND VPWR VPWR VGND clk _01568_ reset_n keymem.key_mem\[4\]\[44\] sky130_fd_sc_hd__dfrtp_2
X_22287_ VGND VPWR _01850_ _06632_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_206_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24026_ VGND VPWR VPWR VGND clk _00519_ reset_n keymem.key_mem\[12\]\[19\] sky130_fd_sc_hd__dfrtp_2
X_12040_ VPWR VGND VPWR VGND _07640_ keymem.key_mem\[9\]\[2\] _07592_ keymem.key_mem\[2\]\[2\]
+ _07546_ _07641_ sky130_fd_sc_hd__a221o_2
XFILLER_0_104_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21238_ VGND VPWR VPWR VGND _06065_ _03434_ keymem.key_mem\[6\]\[92\] _06074_ sky130_fd_sc_hd__mux2_2
XFILLER_0_44_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_178_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21169_ VGND VPWR VPWR VGND _06029_ _03139_ keymem.key_mem\[6\]\[59\] _06038_ sky130_fd_sc_hd__mux2_2
XFILLER_0_244_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_258_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13991_ VPWR VGND VGND VPWR _09463_ _09447_ _09362_ sky130_fd_sc_hd__nand2_2
XFILLER_0_204_106 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_123_2_Right_195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_258_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15730_ VPWR VGND VPWR VGND _11186_ enc_block.block_w0_reg\[23\] _08995_ sky130_fd_sc_hd__or2_2
X_12942_ VGND VPWR enc_block.round_key\[77\] _08467_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24928_ VGND VPWR VPWR VGND clk _01421_ reset_n keymem.key_mem\[5\]\[25\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_1234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_306 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15661_ _10487_ _11118_ _10514_ _10765_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_119_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12873_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[71\] _07711_ keymem.key_mem\[1\]\[71\]
+ _07671_ _08405_ sky130_fd_sc_hd__a22o_2
X_24859_ VGND VPWR VPWR VGND clk _01352_ reset_n keymem.key_mem\[6\]\[84\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_213_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17400_ VPWR VGND VPWR VGND _03484_ _03482_ _03212_ key[227] _03366_ _03485_ sky130_fd_sc_hd__a221o_2
XFILLER_0_51_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14612_ VGND VPWR VGND VPWR _10078_ _10077_ _10079_ _10080_ sky130_fd_sc_hd__a21o_2
XFILLER_0_16_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11824_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[15\] dec_new_block\[79\]
+ _07476_ sky130_fd_sc_hd__mux2_2
X_18380_ VPWR VGND VPWR VGND _04274_ _03970_ _10087_ sky130_fd_sc_hd__or2_2
XFILLER_0_189_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15592_ VGND VPWR keymem.prev_key1_reg\[78\] _11045_ _11050_ _11046_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_115_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17331_ VPWR VGND VGND VPWR _10287_ _03424_ key[219] sky130_fd_sc_hd__nor2_2
X_14543_ VPWR VGND VPWR VGND _10010_ _10011_ _09191_ _09804_ sky130_fd_sc_hd__or3b_2
XFILLER_0_189_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11755_ VGND VPWR result[44] _07441_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_56_748 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_55_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17262_ VPWR VGND key[212] _03362_ _09868_ VPWR VGND sky130_fd_sc_hd__and2_2
X_14474_ VGND VPWR VGND VPWR _09115_ _09217_ _09943_ _09102_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_265_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11686_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[10\] dec_new_block\[10\]
+ _07407_ sky130_fd_sc_hd__mux2_2
X_19001_ VGND VPWR _04831_ enc_block.block_w3_reg\[17\] _04830_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_16213_ VPWR VGND VGND VPWR _11303_ _02378_ _11280_ sky130_fd_sc_hd__nor2_2
XFILLER_0_64_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_265_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13425_ VGND VPWR enc_block.round_key\[125\] _08902_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17193_ VGND VPWR VGND VPWR _11022_ _11021_ _03300_ _03298_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_113_319 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16144_ VPWR VGND VGND VPWR _11219_ _11375_ _11598_ _11386_ _11400_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_140_116 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13356_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[119\] _07743_ keymem.key_mem\[2\]\[119\]
+ _08116_ _08840_ sky130_fd_sc_hd__a22o_2
XFILLER_0_126_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1227 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12307_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[18\] _07535_ _07891_ _07887_ _07892_
+ sky130_fd_sc_hd__o22a_2
X_16075_ VGND VPWR VGND VPWR _11420_ _11296_ _11530_ _11404_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_87_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13287_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[112\] _07659_ keymem.key_mem\[7\]\[112\]
+ _07608_ _08778_ sky130_fd_sc_hd__a22o_2
XFILLER_0_62_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_267_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15026_ VGND VPWR VGND VPWR _10490_ _10483_ _10451_ _10453_ _10464_ sky130_fd_sc_hd__a211o_2
X_19903_ VGND VPWR _00735_ _05363_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12238_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[13\] _07581_ keymem.key_mem\[4\]\[13\]
+ _07550_ _07828_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19834_ VPWR VGND VGND VPWR _05327_ keymem.key_mem\[11\]\[75\] _05243_ sky130_fd_sc_hd__nand2_2
X_12169_ VGND VPWR VGND VPWR _07665_ keymem.key_mem\[4\]\[8\] _07756_ _07758_ _07764_
+ _07763_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_23_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19765_ VGND VPWR VPWR VGND _05281_ keymem.key_mem\[11\]\[42\] _02972_ _05291_ sky130_fd_sc_hd__mux2_2
X_16977_ VGND VPWR VGND VPWR _02682_ _02681_ _03105_ keymem.prev_key1_reg\[56\] sky130_fd_sc_hd__a21oi_2
XFILLER_0_237_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15928_ VPWR VGND VPWR VGND _11265_ _11216_ _11247_ _11166_ _11384_ sky130_fd_sc_hd__or4_2
XFILLER_0_36_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18716_ VPWR VGND VGND VPWR _04512_ _04575_ _04283_ sky130_fd_sc_hd__nor2_2
XFILLER_0_265_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19696_ VGND VPWR VPWR VGND _05247_ keymem.key_mem\[11\]\[9\] _10747_ _05255_ sky130_fd_sc_hd__mux2_2
X_18647_ VPWR VGND VPWR VGND _04513_ _04459_ _04511_ enc_block.block_w1_reg\[21\]
+ _04424_ _00329_ sky130_fd_sc_hd__a221o_2
X_15859_ VGND VPWR VGND VPWR _11311_ _11303_ _11314_ _11308_ _11315_ sky130_fd_sc_hd__o22a_2
XFILLER_0_91_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_531 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_204_695 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_133_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18578_ VGND VPWR VGND VPWR _04450_ _03951_ _04451_ _00322_ sky130_fd_sc_hd__a21o_2
XFILLER_0_52_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_1029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17529_ VPWR VGND VPWR VGND _03596_ key[117] _11543_ sky130_fd_sc_hd__or2_2
XFILLER_0_86_383 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_52_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20540_ VGND VPWR VPWR VGND _05692_ _02607_ keymem.key_mem\[8\]\[22\] _05702_ sky130_fd_sc_hd__mux2_2
XFILLER_0_34_409 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_116_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20471_ VGND VPWR VPWR VGND _05660_ _03607_ keymem.key_mem\[9\]\[118\] _05665_ sky130_fd_sc_hd__mux2_2
XFILLER_0_116_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22210_ VGND VPWR _01813_ _06592_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_15_656 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23190_ VGND VPWR VPWR VGND _06880_ _07082_ keymem.prev_key1_reg\[126\] _07083_ sky130_fd_sc_hd__mux2_2
XFILLER_0_131_138 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_259_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22141_ VGND VPWR VPWR VGND _06554_ _09724_ keymem.key_mem\[2\]\[1\] _06556_ sky130_fd_sc_hd__mux2_2
XFILLER_0_2_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22072_ VGND VPWR _01749_ _06518_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_220_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21023_ VGND VPWR VPWR VGND _05956_ _05073_ keymem.key_mem\[7\]\[119\] _05960_ sky130_fd_sc_hd__mux2_2
XFILLER_0_61_1095 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25831_ VGND VPWR VPWR VGND clk _02324_ reset_n enc_block.block_w3_reg\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_236_1003 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_173_1304 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_241_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25762_ keymem.prev_key1_reg\[78\] clk _02255_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_184_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22974_ VGND VPWR VGND VPWR _06952_ _02960_ _02958_ _02963_ _06951_ sky130_fd_sc_hd__a211o_2
XFILLER_0_93_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24713_ VGND VPWR VPWR VGND clk _01206_ reset_n keymem.key_mem\[7\]\[66\] sky130_fd_sc_hd__dfrtp_2
X_21925_ VGND VPWR VGND VPWR _06440_ keymem.key_mem_we _02787_ _06432_ _01680_ sky130_fd_sc_hd__a31o_2
XFILLER_0_223_982 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_241_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25693_ keymem.prev_key1_reg\[9\] clk _02186_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_210_610 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24644_ VGND VPWR VPWR VGND clk _01137_ reset_n keymem.key_mem\[8\]\[125\] sky130_fd_sc_hd__dfrtp_2
X_21856_ VGND VPWR _01651_ _06400_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_194_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_139_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20807_ VGND VPWR VGND VPWR _05845_ keymem.key_mem_we _11547_ _05838_ _01157_ sky130_fd_sc_hd__a31o_2
XFILLER_0_37_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21787_ VGND VPWR _01618_ _06364_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24575_ VGND VPWR VPWR VGND clk _01068_ reset_n keymem.key_mem\[8\]\[56\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_320 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_342 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23526_ VGND VPWR VPWR VGND clk _00027_ reset_n keymem.key_mem\[14\]\[15\] sky130_fd_sc_hd__dfrtp_2
X_20738_ VGND VPWR VPWR VGND _05805_ _03592_ keymem.key_mem\[8\]\[116\] _05806_ sky130_fd_sc_hd__mux2_2
XFILLER_0_203_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_241 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23457_ VGND VPWR VGND VPWR _07320_ _07319_ _07322_ _07318_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_110_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20669_ VGND VPWR _01095_ _05769_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_208_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13210_ VPWR VGND VPWR VGND _08708_ keymem.key_mem\[13\]\[104\] _07668_ keymem.key_mem\[14\]\[104\]
+ _07666_ _08709_ sky130_fd_sc_hd__a221o_2
X_22408_ VGND VPWR _06696_ _06695_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14190_ VPWR VGND VPWR VGND _09650_ _09660_ _09654_ _09644_ _09661_ sky130_fd_sc_hd__or4_2
X_23388_ VPWR VGND VPWR VGND _07260_ block[18] _04139_ enc_block.block_w0_reg\[18\]
+ _04138_ _07261_ sky130_fd_sc_hd__a221o_2
XFILLER_0_184_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25127_ VGND VPWR VPWR VGND clk _01620_ reset_n keymem.key_mem\[4\]\[96\] sky130_fd_sc_hd__dfrtp_2
X_13141_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[97\] _08391_ keymem.key_mem\[2\]\[97\]
+ _07646_ _08647_ sky130_fd_sc_hd__a22o_2
X_22339_ VGND VPWR VPWR VGND _06658_ _03459_ keymem.key_mem\[2\]\[95\] _06660_ sky130_fd_sc_hd__mux2_2
XFILLER_0_108_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13072_ VGND VPWR VGND VPWR _08585_ _07839_ keymem.key_mem\[11\]\[90\] _08582_ _08584_
+ sky130_fd_sc_hd__a211o_2
X_25058_ VGND VPWR VPWR VGND clk _01551_ reset_n keymem.key_mem\[4\]\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_130_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16900_ VGND VPWR VPWR VGND _02986_ keymem.key_mem\[14\]\[48\] _03035_ _03036_ sky130_fd_sc_hd__mux2_2
X_12023_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[1\] _07582_ keymem.key_mem\[1\]\[1\]
+ _07624_ _07625_ sky130_fd_sc_hd__a22o_2
X_24009_ VGND VPWR VPWR VGND clk _00502_ reset_n keymem.key_mem\[12\]\[2\] sky130_fd_sc_hd__dfrtp_2
X_17880_ VGND VPWR _03372_ _02484_ _03850_ _03789_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_217_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_79_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16831_ VGND VPWR VPWR VGND _02884_ keymem.key_mem\[14\]\[42\] _02972_ _02973_ sky130_fd_sc_hd__mux2_2
XFILLER_0_79_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1223 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_137_1_Left_404 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_189_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19550_ VGND VPWR VGND VPWR _05176_ keymem.key_mem_we _03235_ _05164_ _00569_ sky130_fd_sc_hd__a31o_2
XFILLER_0_232_223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16762_ VGND VPWR VGND VPWR _09866_ key[164] _02910_ _02909_ sky130_fd_sc_hd__a21oi_2
X_13974_ VGND VPWR VGND VPWR _09446_ _09444_ _09388_ _09441_ _09336_ _09445_ sky130_fd_sc_hd__o221ai_2
X_18501_ VGND VPWR _04382_ _03965_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_124_2_Right_196 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_1031 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15713_ VGND VPWR VGND VPWR _11169_ enc_block.sword_ctr_reg\[0\] enc_block.block_w1_reg\[19\]
+ enc_block.sword_ctr_reg\[1\] sky130_fd_sc_hd__and3b_2
XFILLER_0_191_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19481_ VPWR VGND keymem.key_mem\[12\]\[37\] _05140_ _05128_ VPWR VGND sky130_fd_sc_hd__and2_2
X_12925_ VPWR VGND VPWR VGND _08451_ keymem.key_mem\[6\]\[76\] _07739_ keymem.key_mem\[10\]\[76\]
+ _07865_ _08452_ sky130_fd_sc_hd__a221o_2
XFILLER_0_198_650 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_244_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16693_ VGND VPWR VGND VPWR _02845_ _10360_ _02843_ _02844_ _02846_ sky130_fd_sc_hd__a31o_2
XFILLER_0_87_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18432_ VGND VPWR _04319_ enc_block.block_w2_reg\[17\] enc_block.block_w1_reg\[25\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15644_ VPWR VGND _11101_ keymem.prev_key1_reg\[47\] keymem.prev_key1_reg\[15\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
X_12856_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[69\] _08090_ keymem.key_mem\[1\]\[69\]
+ _07969_ _08390_ sky130_fd_sc_hd__a22o_2
XFILLER_0_87_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_150_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11807_ VGND VPWR result[70] _07467_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_29_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18363_ VPWR VGND VGND VPWR _04258_ _04004_ _09924_ sky130_fd_sc_hd__nand2_2
X_15575_ VPWR VGND VGND VPWR _11034_ _11032_ _11033_ sky130_fd_sc_hd__nand2_2
XFILLER_0_16_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_320 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12787_ VPWR VGND VPWR VGND _08327_ keymem.key_mem\[9\]\[62\] _07919_ keymem.key_mem\[12\]\[62\]
+ _07807_ _08328_ sky130_fd_sc_hd__a221o_2
XFILLER_0_260_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17314_ VPWR VGND VPWR VGND _03408_ _10902_ _03406_ key[217] _03366_ _03409_ sky130_fd_sc_hd__a221o_2
X_14526_ VPWR VGND VGND VPWR _09167_ _09095_ _09994_ _09658_ _09168_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_16_409 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18294_ VPWR VGND VPWR VGND _04196_ _04194_ _04195_ sky130_fd_sc_hd__or2_2
X_11738_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[4\] dec_new_block\[36\]
+ _07433_ sky130_fd_sc_hd__mux2_2
XFILLER_0_113_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_25_910 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_260_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17245_ VGND VPWR _03347_ _03346_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14457_ VPWR VGND VGND VPWR _09926_ keymem.prev_key1_reg\[67\] _09925_ sky130_fd_sc_hd__nand2_2
X_11669_ VGND VPWR result[1] _07398_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_226_1205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_189_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13408_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[124\] _07963_ keymem.key_mem\[8\]\[124\]
+ _07958_ _08887_ sky130_fd_sc_hd__a22o_2
X_17176_ VGND VPWR VPWR VGND _03283_ _02947_ _03285_ _10902_ _03284_ sky130_fd_sc_hd__o211a_2
X_14388_ VPWR VGND VGND VPWR _09854_ _09858_ _09853_ sky130_fd_sc_hd__nor2_2
X_16127_ VGND VPWR VGND VPWR _11270_ _11473_ _11211_ _11320_ _11581_ sky130_fd_sc_hd__o22a_2
XFILLER_0_40_946 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13339_ VGND VPWR VGND VPWR _08016_ keymem.key_mem\[7\]\[117\] _08822_ _08824_ _08825_
+ _08736_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_11_147 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16058_ VPWR VGND VGND VPWR _11235_ _11327_ _11513_ _11219_ _11469_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_267_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15009_ VGND VPWR _10473_ _10397_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_69_1_Left_336 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_97_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19817_ VGND VPWR _00694_ _05318_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_237_1301 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_208_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_58_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_1_Left_388 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_237_1345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_159_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19748_ VGND VPWR _00661_ _05282_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_251_576 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_170_1_Right_771 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19679_ VGND VPWR _00629_ _05245_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_154_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_176_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21710_ VGND VPWR _01581_ _06324_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_52_1017 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22690_ VGND VPWR VPWR VGND _06809_ keymem.key_mem\[0\]\[34\] _02894_ _06816_ sky130_fd_sc_hd__mux2_2
XFILLER_0_154_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_176_344 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21641_ VGND VPWR _01548_ _06288_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_183_1_Left_450 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_74_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_19_247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_69_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24360_ VGND VPWR VPWR VGND clk _00853_ reset_n keymem.key_mem\[10\]\[97\] sky130_fd_sc_hd__dfrtp_2
X_21572_ VGND VPWR _01517_ _06250_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_578 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_151_2_Left_622 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_248_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23311_ VGND VPWR _07192_ _07092_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20523_ VGND VPWR _01025_ _05693_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_69_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24291_ VGND VPWR VPWR VGND clk _00784_ reset_n keymem.key_mem\[10\]\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_248_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23242_ VGND VPWR _07129_ enc_block.block_w3_reg\[31\] enc_block.block_w1_reg\[12\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20454_ VGND VPWR VPWR VGND _05649_ _03555_ keymem.key_mem\[9\]\[110\] _05656_ sky130_fd_sc_hd__mux2_2
XFILLER_0_209_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23173_ VGND VPWR VGND VPWR _03616_ _03615_ _03619_ _07072_ sky130_fd_sc_hd__a21o_2
XFILLER_0_127_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20385_ VGND VPWR VPWR VGND _05614_ _03306_ keymem.key_mem\[9\]\[77\] _05620_ sky130_fd_sc_hd__mux2_2
XFILLER_0_3_870 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_242_1051 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_105_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22124_ VGND VPWR _01774_ _06545_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_88_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_30_489 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_203_1057 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22055_ VGND VPWR _01741_ _06509_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_179_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_377 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21006_ VGND VPWR VPWR VGND _05945_ _05056_ keymem.key_mem\[7\]\[111\] _05951_ sky130_fd_sc_hd__mux2_2
XFILLER_0_255_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_199_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25814_ VGND VPWR VPWR VGND clk _02307_ reset_n enc_block.block_w3_reg\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_216_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25745_ keymem.prev_key1_reg\[61\] clk _02238_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_69_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22957_ VGND VPWR VGND VPWR _02211_ _06941_ _06916_ keymem.prev_key1_reg\[34\] sky130_fd_sc_hd__o21a_2
XFILLER_0_214_1120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12710_ VGND VPWR enc_block.round_key\[54\] _08258_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_167_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21908_ VPWR VGND keymem.key_mem\[3\]\[21\] _06431_ _06427_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13690_ VGND VPWR VPWR VGND _09085_ _09082_ _09105_ _09162_ sky130_fd_sc_hd__or3_2
X_25676_ VGND VPWR VPWR VGND clk _02169_ reset_n keymem.rcon_logic.tmp_rcon\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_116_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22888_ VGND VPWR VPWR VGND _06878_ _06898_ keymem.prev_key1_reg\[8\] _06899_ sky130_fd_sc_hd__mux2_2
X_12641_ VGND VPWR VGND VPWR _07778_ keymem.key_mem\[3\]\[48\] _08192_ _08195_ _08196_
+ _08069_ sky130_fd_sc_hd__a2111o_2
X_24627_ VGND VPWR VPWR VGND clk _01120_ reset_n keymem.key_mem\[8\]\[108\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_194_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21839_ VGND VPWR VPWR VGND _06388_ _03613_ keymem.key_mem\[4\]\[119\] _06392_ sky130_fd_sc_hd__mux2_2
XFILLER_0_13_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_2_Left_554 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15360_ VPWR VGND VGND VPWR _10821_ _10822_ _10820_ sky130_fd_sc_hd__nor2_2
X_12572_ VGND VPWR VGND VPWR _08134_ _08050_ keymem.key_mem\[7\]\[41\] _08130_ _08133_
+ sky130_fd_sc_hd__a211o_2
X_24558_ VGND VPWR VPWR VGND clk _01051_ reset_n keymem.key_mem\[8\]\[39\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14311_ VGND VPWR VGND VPWR _09553_ _09780_ _09372_ _09397_ _09781_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_19_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_266_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23509_ VGND VPWR VPWR VGND clk _00005_ reset_n aes_core_ctrl_reg\[1\] sky130_fd_sc_hd__dfrtp_2
X_15291_ VPWR VGND VGND VPWR _10554_ _10753_ _10513_ sky130_fd_sc_hd__nor2_2
X_24489_ VGND VPWR VPWR VGND clk _00982_ reset_n keymem.key_mem\[9\]\[98\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_184_1230 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_1257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_80_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17030_ VPWR VGND _03153_ _02794_ _02793_ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_11_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14242_ VGND VPWR VGND VPWR _09712_ _09713_ _09711_ _09710_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_80_378 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14173_ VPWR VGND VPWR VGND _09642_ _09643_ _09644_ _09640_ _09641_ sky130_fd_sc_hd__or4b_2
XFILLER_0_68_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13124_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[95\] _08577_ _08631_ _08627_ _08632_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_249_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_162_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18981_ VPWR VGND VGND VPWR _04778_ _04814_ _04232_ sky130_fd_sc_hd__nor2_2
XFILLER_0_81_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17932_ VGND VPWR VPWR VGND _03874_ _03885_ keymem.prev_key0_reg\[101\] _03886_ sky130_fd_sc_hd__mux2_2
X_13055_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[89\] _07656_ keymem.key_mem\[1\]\[89\]
+ _07624_ _08569_ sky130_fd_sc_hd__a22o_2
X_12006_ VGND VPWR _07608_ _07567_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17863_ VGND VPWR VPWR VGND _03836_ _03838_ keymem.prev_key0_reg\[79\] _03839_ sky130_fd_sc_hd__mux2_2
XFILLER_0_79_1153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_121_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19602_ VGND VPWR _00594_ _05203_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_206_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16814_ VPWR VGND _02957_ _10730_ keymem.prev_key0_reg\[105\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_17794_ VPWR VGND VPWR VGND _03116_ _03791_ keymem.prev_key0_reg\[57\] _03788_ _00198_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_92_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19533_ VGND VPWR VGND VPWR _05167_ keymem.key_mem_we _03162_ _05164_ _00561_ sky130_fd_sc_hd__a31o_2
X_16745_ VGND VPWR VPWR VGND _02884_ keymem.key_mem\[14\]\[34\] _02894_ _02895_ sky130_fd_sc_hd__mux2_2
X_13957_ VGND VPWR VGND VPWR _09346_ _09429_ _09414_ _09428_ _09394_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_152_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1097 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_125_2_Right_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_92_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19464_ VGND VPWR VGND VPWR _05130_ keymem.key_mem_we _02812_ _05121_ _00529_ sky130_fd_sc_hd__a31o_2
X_12908_ VPWR VGND VPWR VGND _08436_ keymem.key_mem\[11\]\[74\] _08011_ keymem.key_mem\[10\]\[74\]
+ _07743_ _08437_ sky130_fd_sc_hd__a221o_2
XFILLER_0_48_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16676_ VPWR VGND VPWR VGND _02830_ keymem.prev_key1_reg\[94\] sky130_fd_sc_hd__inv_2
X_13888_ VPWR VGND VGND VPWR _09304_ _09360_ _09303_ sky130_fd_sc_hd__nor2_2
XFILLER_0_5_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15627_ VPWR VGND VGND VPWR _10708_ _11082_ _11083_ _11084_ _11085_ sky130_fd_sc_hd__and4b_2
X_18415_ _08948_ _04304_ enc_block.sword_ctr_reg\[0\] _03972_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__and3_2
X_12839_ VGND VPWR VGND VPWR _08375_ _07800_ keymem.key_mem\[1\]\[67\] _08372_ _08374_
+ sky130_fd_sc_hd__a211o_2
X_19395_ VPWR VGND VGND VPWR _08925_ _05091_ _09538_ sky130_fd_sc_hd__nor2_2
XFILLER_0_201_484 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_118_219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_201_495 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18346_ VPWR VGND VGND VPWR _04243_ _04162_ _04242_ sky130_fd_sc_hd__nand2_2
XFILLER_0_228_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15558_ VGND VPWR VPWR VGND _11015_ _11016_ _11012_ _11017_ sky130_fd_sc_hd__or3_2
X_14509_ VGND VPWR VGND VPWR _09116_ _09658_ _09167_ _09978_ sky130_fd_sc_hd__a21o_2
X_18277_ VPWR VGND VPWR VGND _04180_ _04040_ _04178_ enc_block.block_w0_reg\[18\]
+ _04097_ _00292_ sky130_fd_sc_hd__a221o_2
X_15489_ VGND VPWR VGND VPWR _10530_ _10566_ _10476_ _10593_ _10949_ sky130_fd_sc_hd__o22a_2
XFILLER_0_16_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17228_ VGND VPWR _00092_ _03331_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_163_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_140_77 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_4_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17159_ VGND VPWR _00085_ _03269_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_3_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20170_ VGND VPWR _00860_ _05505_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_126_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_235_Right_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_100_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23860_ VGND VPWR VPWR VGND clk _00353_ reset_n enc_block.block_w2_reg\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_174_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22811_ VGND VPWR _06859_ _03733_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23791_ VGND VPWR VPWR VGND clk _00284_ reset_n enc_block.block_w0_reg\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_170_1307 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_174_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_171_1_Right_772 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_71_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25530_ VGND VPWR VPWR VGND clk _02023_ reset_n keymem.key_mem\[1\]\[115\] sky130_fd_sc_hd__dfrtp_2
X_22742_ VGND VPWR _06836_ _03733_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_71_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25461_ VGND VPWR VPWR VGND clk _01954_ reset_n keymem.key_mem\[1\]\[46\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_176_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_220_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22673_ VGND VPWR VPWR VGND _06798_ keymem.key_mem\[0\]\[25\] _02721_ _06808_ sky130_fd_sc_hd__mux2_2
X_24412_ VGND VPWR VPWR VGND clk _00905_ reset_n keymem.key_mem\[9\]\[21\] sky130_fd_sc_hd__dfrtp_2
X_21624_ VGND VPWR _01540_ _06279_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25392_ VGND VPWR VPWR VGND clk _01885_ reset_n keymem.key_mem\[2\]\[105\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_69_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_973 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_111_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24343_ VGND VPWR VPWR VGND clk _00836_ reset_n keymem.key_mem\[10\]\[80\] sky130_fd_sc_hd__dfrtp_2
X_21555_ VGND VPWR _01509_ _06241_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_63_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20506_ VGND VPWR _01017_ _05684_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21486_ VGND VPWR _01476_ _06205_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24274_ VGND VPWR VPWR VGND clk _00767_ reset_n keymem.key_mem\[10\]\[11\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_185_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23225_ VGND VPWR VGND VPWR _07113_ _04266_ _07095_ _07114_ enc_block.block_w3_reg\[2\]
+ sky130_fd_sc_hd__o2bb2a_2
X_20437_ VGND VPWR VPWR VGND _05638_ _03506_ keymem.key_mem\[9\]\[102\] _05647_ sky130_fd_sc_hd__mux2_2
XFILLER_0_181_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23156_ VGND VPWR VGND VPWR _02289_ _07062_ _06888_ keymem.prev_key1_reg\[112\] sky130_fd_sc_hd__o21a_2
X_20368_ VGND VPWR VPWR VGND _05602_ _03235_ keymem.key_mem\[9\]\[69\] _05611_ sky130_fd_sc_hd__mux2_2
XFILLER_0_261_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_100_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_222_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22107_ VGND VPWR _01766_ _06536_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23087_ VPWR VGND VGND VPWR _07019_ _02653_ _06976_ sky130_fd_sc_hd__nand2_2
XFILLER_0_246_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_235_808 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20299_ VGND VPWR VPWR VGND _05569_ _02913_ keymem.key_mem\[9\]\[36\] _05575_ sky130_fd_sc_hd__mux2_2
X_22038_ VGND VPWR VPWR VGND _06494_ _05002_ keymem.key_mem\[3\]\[81\] _06501_ sky130_fd_sc_hd__mux2_2
XFILLER_0_209_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14860_ VGND VPWR _10325_ _09522_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_192_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13811_ VGND VPWR VGND VPWR enc_block.block_w1_reg\[29\] _08948_ _09022_ _09281_
+ _09283_ _09282_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_243_885 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_216_1226 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14791_ VGND VPWR VGND VPWR _09418_ _09352_ _09495_ _10257_ sky130_fd_sc_hd__a21o_2
X_23989_ VGND VPWR VPWR VGND clk _00482_ reset_n keymem.key_mem\[13\]\[110\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_153_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16530_ VGND VPWR VPWR VGND _02662_ keymem.key_mem\[14\]\[24\] _02689_ _02690_ sky130_fd_sc_hd__mux2_2
X_13742_ VGND VPWR VPWR VGND _09206_ _09213_ _09198_ _09214_ sky130_fd_sc_hd__or3_2
X_25728_ keymem.prev_key1_reg\[44\] clk _02221_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_167_130 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16461_ VGND VPWR VGND VPWR _11352_ _11305_ _11182_ _11399_ _02622_ sky130_fd_sc_hd__o22a_2
X_13673_ VGND VPWR _09145_ _09144_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25659_ VGND VPWR VPWR VGND clk _02152_ reset_n keymem.key_mem\[0\]\[116\] sky130_fd_sc_hd__dfrtp_2
X_18200_ VPWR VGND _04110_ enc_block.block_w2_reg\[15\] enc_block.block_w2_reg\[11\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_6_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15412_ VGND VPWR VPWR VGND _10871_ _10872_ _10870_ _10873_ sky130_fd_sc_hd__or3_2
XFILLER_0_39_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12624_ VGND VPWR VGND VPWR _08181_ _08008_ keymem.key_mem\[2\]\[46\] _08180_ _07896_
+ sky130_fd_sc_hd__a211o_2
X_19180_ VGND VPWR _00421_ _04954_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16392_ VGND VPWR VGND VPWR _11367_ _11311_ _02554_ _11404_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_182_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18131_ VPWR VGND VGND VPWR _04047_ _04044_ _04046_ sky130_fd_sc_hd__nand2_2
X_15343_ VGND VPWR VGND VPWR _10547_ _10513_ _10805_ _10522_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_249_1057 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12555_ VPWR VGND VPWR VGND _08117_ keymem.key_mem\[10\]\[40\] _07786_ keymem.key_mem\[4\]\[40\]
+ _07552_ _08118_ sky130_fd_sc_hd__a221o_2
XFILLER_0_53_356 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18062_ VPWR VGND _03983_ enc_block.block_w3_reg\[7\] enc_block.block_w3_reg\[0\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_0_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15274_ VGND VPWR VGND VPWR _09708_ _09679_ _10737_ keymem.prev_key1_reg\[105\] sky130_fd_sc_hd__a21oi_2
X_12486_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[33\] _07893_ _08055_ _08049_ _08056_
+ sky130_fd_sc_hd__o22a_2
X_17013_ VPWR VGND VPWR VGND _03138_ _10325_ _03135_ _03136_ _03137_ _10281_ sky130_fd_sc_hd__o311a_2
X_14225_ VGND VPWR VGND VPWR _09671_ _09061_ _09693_ _09694_ _09696_ _09695_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_262_1257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_80_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_776 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14156_ VPWR VGND VPWR VGND _09624_ _09626_ _09625_ _09621_ _09627_ sky130_fd_sc_hd__or4_2
XFILLER_0_240_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13107_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[94\] _07716_ keymem.key_mem\[1\]\[94\]
+ _07624_ _08616_ sky130_fd_sc_hd__a22o_2
XFILLER_0_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_240_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14087_ VGND VPWR VGND VPWR _09422_ _09444_ _09391_ _09426_ _09248_ _09558_ sky130_fd_sc_hd__o32a_2
X_18964_ VGND VPWR _04798_ _03952_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_226_808 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17915_ VGND VPWR _03874_ _03673_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13038_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[87\] _08216_ keymem.key_mem\[4\]\[87\]
+ _08077_ _08554_ sky130_fd_sc_hd__a22o_2
XFILLER_0_256_1017 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18895_ VGND VPWR _04736_ enc_block.block_w0_reg\[14\] _04668_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17846_ VGND VPWR VGND VPWR _03274_ keymem.prev_key1_reg\[74\] _03827_ _03818_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_261_660 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_234_1326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_206_598 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14989_ VGND VPWR _10453_ _10452_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17777_ VGND VPWR VPWR VGND _03777_ _03072_ keymem.prev_key0_reg\[52\] _03780_ sky130_fd_sc_hd__mux2_2
XFILLER_0_135_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_233_384 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_88_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_44_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19516_ VGND VPWR _05158_ _05094_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_156_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16728_ VPWR VGND VPWR VGND _02879_ keymem.prev_key1_reg\[33\] sky130_fd_sc_hd__inv_2
XFILLER_0_92_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_126_2_Right_198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_158_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19447_ VGND VPWR _05121_ _05092_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16659_ VGND VPWR _00041_ _02813_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_737 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_201_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_88_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19378_ VGND VPWR VPWR VGND _05067_ _05079_ keymem.key_mem\[13\]\[122\] _05080_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18329_ VGND VPWR _04228_ _04226_ _04227_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_151_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21340_ VGND VPWR _01406_ _06129_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_71_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_464 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21271_ VGND VPWR _01375_ _06091_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_128_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23010_ VGND VPWR _02232_ _06973_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20222_ VGND VPWR _05534_ _05533_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_8_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1285 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_275 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20153_ VGND VPWR _00852_ _05496_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_25_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_616 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_99_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20084_ VGND VPWR _00819_ _05460_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24961_ VGND VPWR VPWR VGND clk _01454_ reset_n keymem.key_mem\[5\]\[58\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_209_370 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23912_ VGND VPWR VPWR VGND clk _00405_ reset_n keymem.key_mem\[13\]\[33\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_88_2_Right_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24892_ VGND VPWR VPWR VGND clk _01385_ reset_n keymem.key_mem\[6\]\[117\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_217_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_885 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23843_ VGND VPWR VPWR VGND clk _00336_ reset_n enc_block.block_w1_reg\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_1089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_135_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_79_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_196_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23774_ VGND VPWR VPWR VGND clk _00000_ reset_n enc_block.enc_ctrl_reg\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_79_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20986_ VGND VPWR _01241_ _05940_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_135_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_172_1_Right_773 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25513_ VGND VPWR VPWR VGND clk _02006_ reset_n keymem.key_mem\[1\]\[98\] sky130_fd_sc_hd__dfrtp_2
X_22725_ VGND VPWR _02093_ _06827_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_71_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_137_303 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25444_ VGND VPWR VPWR VGND clk _01937_ reset_n keymem.key_mem\[1\]\[29\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_164_111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22656_ VGND VPWR _02052_ _06799_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21607_ VGND VPWR _01532_ _06270_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25375_ VGND VPWR VPWR VGND clk _01868_ reset_n keymem.key_mem\[2\]\[88\] sky130_fd_sc_hd__dfrtp_2
X_22587_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[101\] _06767_ _06766_ _05035_ _02009_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_62_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_211_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24326_ VGND VPWR VPWR VGND clk _00819_ reset_n keymem.key_mem\[10\]\[63\] sky130_fd_sc_hd__dfrtp_2
X_12340_ VGND VPWR VGND VPWR _07793_ keymem.key_mem\[0\]\[20\] _07922_ _07916_ _07911_
+ _07923_ sky130_fd_sc_hd__o32a_2
X_21538_ VGND VPWR VPWR VGND _06231_ _03525_ keymem.key_mem\[5\]\[105\] _06233_ sky130_fd_sc_hd__mux2_2
XFILLER_0_211_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_146_1_Left_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_146_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24257_ VGND VPWR VPWR VGND clk _00750_ reset_n keymem.key_mem\[11\]\[122\] sky130_fd_sc_hd__dfrtp_2
X_12271_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[15\] _07645_ _07858_ _07852_ _07859_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_160_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21469_ VGND VPWR VPWR VGND _06196_ _03259_ keymem.key_mem\[5\]\[72\] _06197_ sky130_fd_sc_hd__mux2_2
XFILLER_0_146_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14010_ VPWR VGND VGND VPWR _09357_ _09366_ _09482_ _09434_ _09380_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_31_551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23208_ VPWR VGND _07098_ enc_block.block_w2_reg\[7\] enc_block.block_w2_reg\[0\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_120_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_142_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24188_ VGND VPWR VPWR VGND clk _00681_ reset_n keymem.key_mem\[11\]\[53\] sky130_fd_sc_hd__dfrtp_2
X_23139_ VGND VPWR _02283_ _07051_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_43_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15961_ VGND VPWR VGND VPWR _11417_ _11273_ _11228_ _11227_ _11226_ sky130_fd_sc_hd__and4_2
X_17700_ VGND VPWR _03731_ _03728_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14912_ VGND VPWR VPWR VGND _10373_ _10374_ keymem.prev_key1_reg\[72\] _10376_ sky130_fd_sc_hd__or3_2
X_15892_ VGND VPWR VGND VPWR _11348_ _11258_ _11286_ _11174_ _11263_ sky130_fd_sc_hd__and4_2
X_18680_ VPWR VGND VPWR VGND _04542_ _04459_ _04541_ enc_block.block_w1_reg\[25\]
+ _04328_ _00333_ sky130_fd_sc_hd__a221o_2
XFILLER_0_262_468 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_76_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14843_ VGND VPWR VPWR VGND _10308_ _09303_ _09447_ _09312_ _10307_ sky130_fd_sc_hd__o31a_2
X_17631_ VGND VPWR VGND VPWR _09869_ keymem.prev_key1_reg\[3\] _03683_ _03670_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_243_682 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_157_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_153_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17562_ VPWR VGND VGND VPWR _10287_ _03625_ key[249] sky130_fd_sc_hd__nor2_2
X_14774_ VGND VPWR VGND VPWR _09375_ _09474_ _09552_ _09335_ _09331_ _10240_ sky130_fd_sc_hd__o32a_2
X_11986_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[0\] _07588_ keymem.key_mem\[14\]\[0\]
+ _07584_ _07589_ sky130_fd_sc_hd__a22o_2
XFILLER_0_187_247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_114_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19301_ VGND VPWR VPWR VGND _05025_ _05027_ keymem.key_mem\[13\]\[97\] _05028_ sky130_fd_sc_hd__mux2_2
XFILLER_0_153_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16513_ VGND VPWR _02673_ keymem.prev_key0_reg\[56\] keymem.prev_key0_reg\[88\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13725_ VGND VPWR VGND VPWR _09197_ _09196_ _09105_ _09177_ _09167_ sky130_fd_sc_hd__a211o_2
X_17493_ VGND VPWR VGND VPWR _03565_ _03564_ _03563_ _10092_ sky130_fd_sc_hd__o21a_2
XFILLER_0_6_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16444_ VGND VPWR VGND VPWR keylen _02606_ _02605_ keymem.prev_key1_reg\[22\] _02601_
+ _02603_ sky130_fd_sc_hd__a311oi_2
X_19232_ VPWR VGND keymem.key_mem\[13\]\[71\] _04985_ _04979_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_2_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13656_ VGND VPWR VPWR VGND _09014_ _08991_ _09043_ _09128_ sky130_fd_sc_hd__or3_2
XFILLER_0_6_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19163_ VPWR VGND keymem.key_mem_we _04943_ _02998_ VPWR VGND sky130_fd_sc_hd__and2_2
X_12607_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[45\] _07667_ keymem.key_mem\[4\]\[45\]
+ _07551_ _08165_ sky130_fd_sc_hd__a22o_2
XFILLER_0_2_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16375_ VGND VPWR VPWR VGND _10993_ _11018_ keymem.round_ctr_reg\[0\] _02538_ sky130_fd_sc_hd__or3_2
X_13587_ VPWR VGND VGND VPWR _09058_ _09059_ _09057_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_78_1_Left_345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_143_317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_53_131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18114_ VGND VPWR VGND VPWR _04029_ _03951_ _04031_ _00278_ sky130_fd_sc_hd__a21o_2
X_15326_ VGND VPWR VGND VPWR _10633_ _10504_ _10612_ _10530_ _10788_ sky130_fd_sc_hd__o22a_2
X_12538_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[38\] _07668_ keymem.key_mem\[7\]\[38\]
+ _07703_ _08103_ sky130_fd_sc_hd__a22o_2
X_19094_ VGND VPWR VGND VPWR _04901_ keymem.key_mem_we _11447_ _04896_ _00388_ sky130_fd_sc_hd__a31o_2
XPHY_EDGE_ROW_130_1_Left_397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_164_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18045_ VGND VPWR VGND VPWR _03964_ _03963_ _03967_ _03966_ sky130_fd_sc_hd__a21oi_2
X_15257_ VPWR VGND VPWR VGND _10717_ _10719_ _10720_ _10715_ _10716_ sky130_fd_sc_hd__or4b_2
XFILLER_0_125_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_258_708 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12469_ VGND VPWR VGND VPWR _07968_ keymem.key_mem\[9\]\[32\] _08037_ _08039_ _08040_
+ _07574_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_164_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14208_ VGND VPWR VGND VPWR _09669_ _09678_ _09679_ _09661_ _09677_ sky130_fd_sc_hd__nor4_2
XFILLER_0_257_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_199_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15188_ VGND VPWR VGND VPWR _10617_ _10651_ _10652_ _10582_ _10632_ sky130_fd_sc_hd__nor4_2
XFILLER_0_50_882 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_65_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_125_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14139_ VPWR VGND VPWR VGND _09608_ _09609_ _09610_ _09324_ _09607_ sky130_fd_sc_hd__or4b_2
XFILLER_0_22_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_752 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_199_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19996_ VGND VPWR _00777_ _05414_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18947_ VGND VPWR _04783_ _04711_ _04782_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_160_2_Left_631 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18878_ _04719_ _04721_ _04718_ _04720_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_253_479 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_222_822 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17829_ VGND VPWR _00209_ _03815_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_175_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_490 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_171_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20840_ VGND VPWR VPWR VGND _05820_ _04922_ keymem.key_mem\[7\]\[33\] _05863_ sky130_fd_sc_hd__mux2_2
XFILLER_0_178_236 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_72_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_171_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_127_2_Right_199 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_251_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20771_ VPWR VGND keymem.key_mem\[7\]\[1\] _05826_ _05824_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_71_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22510_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[55\] _06737_ _06736_ _04963_ _01963_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_186_280 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23490_ VGND VPWR _07351_ enc_block.block_w2_reg\[6\] _07350_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_278 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_119_358 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22441_ VGND VPWR VPWR VGND _06702_ keymem.key_mem\[1\]\[15\] _11149_ _06714_ sky130_fd_sc_hd__mux2_2
XFILLER_0_44_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_44_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25160_ VGND VPWR VPWR VGND clk _01653_ reset_n keymem.key_mem\[3\]\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_613 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22372_ VGND VPWR VPWR VGND _06669_ _03560_ keymem.key_mem\[2\]\[111\] _06677_ sky130_fd_sc_hd__mux2_2
XFILLER_0_33_849 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_182_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24111_ VGND VPWR VPWR VGND clk _00604_ reset_n keymem.key_mem\[12\]\[104\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_44_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21323_ VGND VPWR _01398_ _06120_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25091_ VGND VPWR VPWR VGND clk _01584_ reset_n keymem.key_mem\[4\]\[60\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_143_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_182_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24042_ VGND VPWR VPWR VGND clk _00535_ reset_n keymem.key_mem\[12\]\[35\] sky130_fd_sc_hd__dfrtp_2
X_21254_ VGND VPWR _01367_ _06082_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_248_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_143_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20205_ VGND VPWR _00877_ _05523_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_40_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21185_ VGND VPWR _01334_ _06046_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_198_1037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_229_465 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_99_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20136_ VGND VPWR _00844_ _05487_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_92_2_Left_563 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_216_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20067_ VGND VPWR _00811_ _05451_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24944_ VGND VPWR VPWR VGND clk _01437_ reset_n keymem.key_mem\[5\]\[41\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_89_2_Right_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24875_ VGND VPWR VPWR VGND clk _01368_ reset_n keymem.key_mem\[6\]\[100\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_240_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_169_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_139_1190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11840_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[23\] dec_new_block\[87\]
+ _07484_ sky130_fd_sc_hd__mux2_2
X_23826_ VGND VPWR VPWR VGND clk _00319_ reset_n enc_block.block_w1_reg\[11\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_240_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_36_1140 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_150_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23757_ keymem.prev_key0_reg\[113\] clk _00254_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_11771_ VGND VPWR result[52] _07449_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_230_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20969_ VGND VPWR VGND VPWR _05931_ keymem.key_mem_we _03444_ _05916_ _01233_ sky130_fd_sc_hd__a31o_2
XFILLER_0_7_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_173_1_Right_774 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13510_ VGND VPWR VGND VPWR _08982_ _08981_ _08980_ keymem.prev_key1_reg\[6\] _08969_
+ _08964_ sky130_fd_sc_hd__a32o_2
XFILLER_0_184_239 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_32_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22708_ VGND VPWR VPWR VGND _06809_ keymem.key_mem\[0\]\[47\] _03025_ _06821_ sky130_fd_sc_hd__mux2_2
XFILLER_0_230_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14490_ VGND VPWR VGND VPWR _09007_ _09072_ _09115_ _09079_ _09959_ sky130_fd_sc_hd__o22a_2
XFILLER_0_3_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23688_ keymem.prev_key0_reg\[44\] clk _00185_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_36_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_306 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25427_ VGND VPWR VPWR VGND clk _01920_ reset_n keymem.key_mem\[1\]\[12\] sky130_fd_sc_hd__dfrtp_2
X_13441_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[127\] _07565_ keymem.key_mem\[11\]\[127\]
+ _07861_ _08917_ sky130_fd_sc_hd__a22o_2
XFILLER_0_3_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22639_ VGND VPWR VPWR VGND _06785_ keymem.key_mem\[0\]\[8\] _10662_ _06791_ sky130_fd_sc_hd__mux2_2
XFILLER_0_137_199 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16160_ VGND VPWR VGND VPWR _11318_ _11235_ _11325_ _11305_ _11614_ sky130_fd_sc_hd__a31o_2
XFILLER_0_1_1160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25358_ VGND VPWR VPWR VGND clk _01851_ reset_n keymem.key_mem\[2\]\[71\] sky130_fd_sc_hd__dfrtp_2
X_13372_ VPWR VGND VPWR VGND _08854_ keymem.key_mem\[11\]\[120\] _08011_ keymem.key_mem\[1\]\[120\]
+ _07671_ _08855_ sky130_fd_sc_hd__a221o_2
XFILLER_0_24_838 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15111_ VGND VPWR _10575_ _10462_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_140_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24309_ VGND VPWR VPWR VGND clk _00802_ reset_n keymem.key_mem\[10\]\[46\] sky130_fd_sc_hd__dfrtp_2
X_12323_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[19\] _07893_ _07906_ _07897_ _07907_
+ sky130_fd_sc_hd__o22a_2
X_16091_ VPWR VGND VPWR VGND _11545_ _09638_ _11457_ key[145] _11043_ _11546_ sky130_fd_sc_hd__a221o_2
XFILLER_0_133_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25289_ VGND VPWR VPWR VGND clk _01782_ reset_n keymem.key_mem\[2\]\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_267_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15042_ VPWR VGND VPWR VGND _10424_ _10435_ _10429_ _10442_ _10506_ sky130_fd_sc_hd__or4_2
XFILLER_0_50_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12254_ VGND VPWR _07843_ _07601_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_82_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19850_ VGND VPWR _00710_ _05335_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_76_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12185_ VGND VPWR _07778_ _07603_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_43_1166 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_43_1177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18801_ VPWR VGND VPWR VGND _04651_ block[37] _04576_ enc_block.block_w1_reg\[5\]
+ _04543_ _04652_ sky130_fd_sc_hd__a221o_2
XFILLER_0_263_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_402 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_78_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19781_ VGND VPWR _00677_ _05299_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16993_ VGND VPWR VPWR VGND _03084_ keymem.key_mem\[14\]\[57\] _03119_ _03120_ sky130_fd_sc_hd__mux2_2
X_18732_ VPWR VGND _04589_ _04588_ enc_block.round_key\[95\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15944_ VGND VPWR _11400_ _11399_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15875_ VGND VPWR VPWR VGND _11173_ _11247_ _11166_ _11331_ sky130_fd_sc_hd__or3_2
X_18663_ VPWR VGND VGND VPWR _04512_ _04528_ _04232_ sky130_fd_sc_hd__nor2_2
X_14826_ VGND VPWR VGND VPWR _09597_ _10291_ _10289_ _10290_ _09764_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_116_46 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_203_343 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17614_ VGND VPWR VGND VPWR _07369_ ready _00140_ _07370_ sky130_fd_sc_hd__a21bo_2
X_18594_ VPWR VGND VPWR VGND _04465_ block[80] _03958_ enc_block.block_w2_reg\[16\]
+ _03953_ _04466_ sky130_fd_sc_hd__a221o_2
XFILLER_0_118_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14757_ VPWR VGND VGND VPWR _09114_ _10223_ _09091_ sky130_fd_sc_hd__nor2_2
X_17545_ VPWR VGND VGND VPWR _03610_ _02651_ _02652_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11969_ VGND VPWR _07572_ _07571_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_175_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_779 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13708_ VPWR VGND VGND VPWR _09033_ _09180_ _09156_ sky130_fd_sc_hd__nor2_2
XFILLER_0_132_12 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_280 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17476_ VGND VPWR VPWR VGND _03534_ keymem.key_mem\[14\]\[109\] _03550_ _03551_ sky130_fd_sc_hd__mux2_2
X_14688_ VGND VPWR VGND VPWR _09012_ _09228_ _10152_ _10153_ _10155_ _10154_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_6_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19215_ VGND VPWR VGND VPWR _04974_ keymem.key_mem_we _03194_ _04968_ _00436_ sky130_fd_sc_hd__a31o_2
X_13639_ VGND VPWR VGND VPWR _09109_ _09033_ _09019_ _09110_ _09111_ sky130_fd_sc_hd__o22a_2
X_16427_ VGND VPWR VPWR VGND keymem.prev_key0_reg\[118\] _02587_ _02589_ _02552_ sky130_fd_sc_hd__a21boi_2
XPHY_EDGE_ROW_17_Left_285 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_116_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_985 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16358_ VGND VPWR VGND VPWR _11316_ _11303_ _11211_ _11320_ _02521_ sky130_fd_sc_hd__o22a_2
X_19146_ VGND VPWR VPWR VGND _04928_ _04931_ keymem.key_mem\[13\]\[38\] _04932_ sky130_fd_sc_hd__mux2_2
XFILLER_0_26_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15309_ VPWR VGND VPWR VGND _10771_ _10443_ _10457_ _10435_ _10609_ _10508_ sky130_fd_sc_hd__o311a_2
XFILLER_0_81_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16289_ VGND VPWR VGND VPWR _11314_ _11327_ _11466_ _11330_ _02453_ sky130_fd_sc_hd__o22a_2
X_19077_ VPWR VGND keymem.key_mem\[13\]\[9\] _04892_ _04887_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_42_679 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_125_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18028_ VGND VPWR _03950_ _03949_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_164_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_521 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_65_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1335 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_160_1158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_275 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_22_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19979_ VGND VPWR _00769_ _05405_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_26_Left_294 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_201_1177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_254_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22990_ VGND VPWR VGND VPWR _06962_ _03019_ _03860_ _06924_ _03023_ sky130_fd_sc_hd__a211o_2
X_21941_ VGND VPWR _06449_ _06402_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_222_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_173_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24660_ VGND VPWR VPWR VGND clk _01153_ reset_n keymem.key_mem\[7\]\[13\] sky130_fd_sc_hd__dfrtp_2
X_21872_ VGND VPWR VGND VPWR _06411_ keymem.key_mem_we _10099_ _06404_ _01656_ sky130_fd_sc_hd__a31o_2
XFILLER_0_136_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23611_ VGND VPWR VPWR VGND clk _00112_ reset_n keymem.key_mem\[14\]\[100\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_72_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20823_ VPWR VGND keymem.key_mem\[7\]\[25\] _05854_ _05844_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_210_847 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24591_ VGND VPWR VPWR VGND clk _01084_ reset_n keymem.key_mem\[8\]\[72\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_106_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23542_ VGND VPWR VPWR VGND clk _00043_ reset_n keymem.key_mem\[14\]\[31\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20754_ VGND VPWR VPWR VGND _05805_ _03647_ keymem.key_mem\[8\]\[124\] _05814_ sky130_fd_sc_hd__mux2_2
X_23473_ VGND VPWR _07336_ _07274_ _07335_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20685_ VGND VPWR VPWR VGND _05772_ _03426_ keymem.key_mem\[8\]\[91\] _05778_ sky130_fd_sc_hd__mux2_2
X_25212_ VGND VPWR VPWR VGND clk _01705_ reset_n keymem.key_mem\[3\]\[53\] sky130_fd_sc_hd__dfrtp_2
X_22424_ VGND VPWR _01914_ _06705_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_33_624 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_169_1194 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_60_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25143_ VGND VPWR VPWR VGND clk _01636_ reset_n keymem.key_mem\[4\]\[112\] sky130_fd_sc_hd__dfrtp_2
X_22355_ VGND VPWR VPWR VGND _06658_ _03511_ keymem.key_mem\[2\]\[103\] _06668_ sky130_fd_sc_hd__mux2_2
XFILLER_0_206_1033 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_108_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21306_ VGND VPWR _01392_ _06109_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_143_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25074_ VGND VPWR VPWR VGND clk _01567_ reset_n keymem.key_mem\[4\]\[43\] sky130_fd_sc_hd__dfrtp_2
X_22286_ VGND VPWR VPWR VGND _06622_ _03245_ keymem.key_mem\[2\]\[70\] _06632_ sky130_fd_sc_hd__mux2_2
XFILLER_0_104_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1077 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_44_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24025_ VGND VPWR VPWR VGND clk _00518_ reset_n keymem.key_mem\[12\]\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_143_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21237_ VGND VPWR _01359_ _06073_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_40_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_217_402 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_44_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21168_ VGND VPWR _01326_ _06037_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_257_593 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_258_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_79_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20119_ VGND VPWR _00836_ _05478_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13990_ VPWR VGND VPWR VGND _09459_ _09461_ _09460_ _09458_ _09462_ sky130_fd_sc_hd__or4_2
XFILLER_0_258_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21099_ VGND VPWR _01293_ _06001_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_77_1251 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12941_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[77\] _08124_ _08466_ _08462_ _08467_
+ sky130_fd_sc_hd__o22a_2
X_24927_ VGND VPWR VPWR VGND clk _01420_ reset_n keymem.key_mem\[5\]\[24\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_99_145 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_225_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_843 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15660_ VGND VPWR VGND VPWR _10527_ _10619_ _11117_ _10628_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_38_1246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24858_ VGND VPWR VPWR VGND clk _01351_ reset_n keymem.key_mem\[6\]\[83\] sky130_fd_sc_hd__dfrtp_2
X_12872_ VGND VPWR enc_block.round_key\[70\] _08404_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_197_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_115_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_197_353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14611_ VPWR VGND _10079_ keymem.prev_key0_reg\[68\] keymem.prev_key0_reg\[36\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
X_11823_ VGND VPWR result[78] _07475_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23809_ VGND VPWR VPWR VGND clk _00302_ reset_n enc_block.block_w0_reg\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_90_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15591_ VPWR VGND _11049_ keymem.prev_key1_reg\[46\] keymem.prev_key1_reg\[14\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_115_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1086 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24789_ VGND VPWR VPWR VGND clk _01282_ reset_n keymem.key_mem\[6\]\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_189_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17330_ VGND VPWR VGND VPWR _02758_ _02757_ _03423_ _02708_ sky130_fd_sc_hd__a21oi_2
X_14542_ VGND VPWR VGND VPWR _09097_ _09079_ _09077_ _09011_ _09230_ _10010_ sky130_fd_sc_hd__o32a_2
X_11754_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[12\] dec_new_block\[44\]
+ _07441_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_51_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_174_1_Right_775 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17261_ VGND VPWR VPWR VGND _03361_ _10735_ _03358_ _03359_ _03360_ sky130_fd_sc_hd__o31a_2
X_14473_ VGND VPWR VGND VPWR _09209_ _08972_ _09942_ _09121_ sky130_fd_sc_hd__a21oi_2
X_11685_ VGND VPWR result[9] _07406_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_265_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16212_ VPWR VGND VPWR VGND _02376_ _02377_ _02374_ _02375_ sky130_fd_sc_hd__or3b_2
X_19000_ VGND VPWR _04830_ enc_block.block_w3_reg\[18\] enc_block.block_w1_reg\[2\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_187_1261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13424_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[125\] _08027_ _08901_ _08897_ _08902_
+ sky130_fd_sc_hd__o22a_2
X_17192_ _11021_ _03299_ _03298_ _11022_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_265_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_63_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16143_ VPWR VGND VGND VPWR _11253_ _11219_ _11597_ _11306_ _11379_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13355_ VGND VPWR enc_block.round_key\[118\] _08839_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_183_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_11_307 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_133_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12306_ VGND VPWR VGND VPWR _07891_ _07547_ keymem.key_mem\[2\]\[18\] _07888_ _07890_
+ sky130_fd_sc_hd__a211o_2
X_16074_ VGND VPWR VGND VPWR _11316_ _11245_ _11529_ _11204_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_1397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_126_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13286_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[112\] _07652_ keymem.key_mem\[14\]\[112\]
+ _08003_ _08777_ sky130_fd_sc_hd__a22o_2
XFILLER_0_122_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15025_ VGND VPWR _10489_ _10488_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19902_ VGND VPWR VPWR VGND _05361_ keymem.key_mem\[11\]\[107\] _03538_ _05363_ sky130_fd_sc_hd__mux2_2
XFILLER_0_62_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12237_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[13\] _07599_ keymem.key_mem\[12\]\[13\]
+ _07620_ _07827_ sky130_fd_sc_hd__a22o_2
XFILLER_0_202_1420 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_23_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19833_ VGND VPWR _05326_ _03279_ _00702_ _05243_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_202_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12168_ VPWR VGND VPWR VGND _07762_ keymem.key_mem\[6\]\[8\] _07760_ keymem.key_mem\[2\]\[8\]
+ _07547_ _07763_ sky130_fd_sc_hd__a221o_2
XFILLER_0_237_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_202_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19764_ VGND VPWR _00669_ _05290_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_236_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12099_ VGND VPWR _07697_ _07545_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16976_ _02681_ _03104_ keymem.prev_key1_reg\[56\] _02682_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_18715_ VPWR VGND _04574_ _04573_ enc_block.round_key\[93\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_237_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15927_ VPWR VGND VPWR VGND _11383_ _11374_ _11382_ sky130_fd_sc_hd__or2_2
XFILLER_0_223_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19695_ VGND VPWR _00636_ _05254_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_36_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18646_ VPWR VGND VGND VPWR _04512_ _04513_ _04211_ sky130_fd_sc_hd__nor2_2
XFILLER_0_258_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15858_ VGND VPWR _11314_ _11313_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_133_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1284 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14809_ VGND VPWR keymem.prev_key1_reg\[70\] _10273_ _10275_ _10274_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_18577_ VGND VPWR VPWR VGND _04316_ enc_block.block_w1_reg\[14\] _04135_ _04451_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_133_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15789_ VGND VPWR _11245_ _11244_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_15_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17528_ VGND VPWR VPWR VGND _02539_ _02540_ _09932_ _03595_ sky130_fd_sc_hd__or3_2
XFILLER_0_15_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_930 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_86_395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_163_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_6_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17459_ VGND VPWR _03302_ key[107] _03536_ _11109_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_20470_ VGND VPWR _01001_ _05664_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_89_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_432 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19129_ VGND VPWR VPWR VGND _04877_ _04920_ keymem.key_mem\[13\]\[32\] _04921_ sky130_fd_sc_hd__mux2_2
XFILLER_0_15_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_246_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_259_836 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22140_ VGND VPWR _01780_ _06555_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_30_649 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_207_1386 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_140_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22071_ VGND VPWR VPWR VGND _06516_ _05027_ keymem.key_mem\[3\]\[97\] _06518_ sky130_fd_sc_hd__mux2_2
XFILLER_0_26_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_891 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21022_ VGND VPWR _01258_ _05959_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_220_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25830_ VGND VPWR VPWR VGND clk _02323_ reset_n enc_block.block_w3_reg\[18\] sky130_fd_sc_hd__dfrtp_2
X_25761_ keymem.prev_key1_reg\[77\] clk _02254_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22973_ VGND VPWR _06951_ _06924_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24712_ VGND VPWR VPWR VGND clk _01205_ reset_n keymem.key_mem\[7\]\[65\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_69_318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21924_ VPWR VGND keymem.key_mem\[3\]\[28\] _06440_ _06439_ VPWR VGND sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_155_1_Left_422 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25692_ keymem.prev_key1_reg\[8\] clk _02185_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_214_1313 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_214_1335 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_136_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24643_ VGND VPWR VPWR VGND clk _01136_ reset_n keymem.key_mem\[8\]\[124\] sky130_fd_sc_hd__dfrtp_2
X_21855_ VGND VPWR VPWR VGND _06262_ _03668_ keymem.key_mem\[4\]\[127\] _06400_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_43_Left_311 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20806_ VPWR VGND keymem.key_mem\[7\]\[17\] _05845_ _05844_ VPWR VGND sky130_fd_sc_hd__and2_2
X_24574_ VGND VPWR VPWR VGND clk _01067_ reset_n keymem.key_mem\[8\]\[55\] sky130_fd_sc_hd__dfrtp_2
X_21786_ VGND VPWR VPWR VGND _06355_ _03452_ keymem.key_mem\[4\]\[94\] _06364_ sky130_fd_sc_hd__mux2_2
XFILLER_0_19_930 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_154_209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23525_ VGND VPWR VPWR VGND clk _00026_ reset_n keymem.key_mem\[14\]\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_194_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20737_ VGND VPWR _05805_ _05675_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_14_Right_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_147_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_92_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_147_294 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_52_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23456_ _07319_ _07321_ _07318_ _07320_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_20668_ VGND VPWR VPWR VGND _05761_ _03355_ keymem.key_mem\[8\]\[83\] _05769_ sky130_fd_sc_hd__mux2_2
XFILLER_0_162_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_208_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22407_ VPWR VGND VGND VPWR _06695_ keymem.key_mem_we _02947_ sky130_fd_sc_hd__nand2_2
XFILLER_0_34_977 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23387_ _07258_ _07260_ _04064_ _07259_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_249_Right_118 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20599_ VGND VPWR VPWR VGND _05725_ _03056_ keymem.key_mem\[8\]\[50\] _05733_ sky130_fd_sc_hd__mux2_2
XFILLER_0_34_999 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25126_ VGND VPWR VPWR VGND clk _01619_ reset_n keymem.key_mem\[4\]\[95\] sky130_fd_sc_hd__dfrtp_2
X_13140_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[97\] _07668_ keymem.key_mem\[6\]\[97\]
+ _07818_ _08646_ sky130_fd_sc_hd__a22o_2
X_22338_ VGND VPWR _01874_ _06659_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_638 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_52_Left_320 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_60_284 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13071_ VPWR VGND VPWR VGND _08583_ keymem.key_mem\[5\]\[90\] _08052_ keymem.key_mem\[1\]\[90\]
+ _07671_ _08584_ sky130_fd_sc_hd__a221o_2
X_25057_ VGND VPWR VPWR VGND clk _01550_ reset_n keymem.key_mem\[4\]\[26\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_159 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22269_ VGND VPWR _01841_ _06623_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_44_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24008_ VGND VPWR VPWR VGND clk _00501_ reset_n keymem.key_mem\[12\]\[1\] sky130_fd_sc_hd__dfrtp_2
X_12022_ VGND VPWR _07624_ _07555_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_23_Right_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_178_1227 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_118_2_Left_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_218_766 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_79_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16830_ VPWR VGND VPWR VGND _02971_ _02967_ _02966_ key[170] _02875_ _02972_ sky130_fd_sc_hd__a221o_2
XFILLER_0_205_427 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_79_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13973_ VGND VPWR VGND VPWR _09381_ _09396_ _09404_ _09423_ _09445_ sky130_fd_sc_hd__a31o_2
XPHY_EDGE_ROW_87_1_Left_354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16761_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[68\] keymem.prev_key1_reg\[36\]
+ _02909_ _02908_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_232_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18500_ VPWR VGND VPWR VGND _04381_ _04291_ _04379_ enc_block.block_w1_reg\[6\] _04317_
+ _00314_ sky130_fd_sc_hd__a221o_2
XFILLER_0_189_139 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15712_ enc_block.sword_ctr_reg\[1\] _11168_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[19\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_12924_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[76\] _07806_ keymem.key_mem\[2\]\[76\]
+ _07697_ _08451_ sky130_fd_sc_hd__a22o_2
X_16692_ VGND VPWR VGND VPWR _10315_ _10292_ _02845_ _09240_ sky130_fd_sc_hd__a21oi_2
X_19480_ VGND VPWR _00536_ _05139_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_232_279 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_115_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_780 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18431_ VPWR VGND _04318_ enc_block.block_w0_reg\[7\] enc_block.block_w0_reg\[0\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_119_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12855_ VGND VPWR VGND VPWR _07835_ keymem.key_mem\[13\]\[69\] _08386_ _08388_ _08389_
+ _08243_ sky130_fd_sc_hd__a2111o_2
X_15643_ VGND VPWR _00026_ _11100_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_244_98 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_115_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11806_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[6\] dec_new_block\[70\]
+ _07467_ sky130_fd_sc_hd__mux2_2
X_18362_ VPWR VGND VPWR VGND _04257_ _04189_ _04255_ enc_block.block_w0_reg\[26\]
+ _03993_ _00300_ sky130_fd_sc_hd__a221o_2
X_15574_ VGND VPWR VPWR VGND _11033_ keymem.prev_key1_reg\[77\] _11030_ _11031_ _09729_
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_150_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Right_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12786_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[62\] _07843_ keymem.key_mem\[4\]\[62\]
+ _07913_ _08327_ sky130_fd_sc_hd__a22o_2
XFILLER_0_29_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1509 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_95_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_230_1170 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14525_ VGND VPWR _00015_ _09993_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17313_ VGND VPWR VGND VPWR keylen _03408_ _03407_ _10323_ _02712_ _02713_ sky130_fd_sc_hd__a311oi_2
X_11737_ VGND VPWR result[35] _07432_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18293_ VPWR VGND _04195_ _04110_ enc_block.block_w0_reg\[28\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_56_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_175_1_Right_776 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_760 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14456_ VPWR VGND _09925_ _09924_ keymem.prev_key1_reg\[99\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_17244_ VGND VPWR VGND VPWR _03346_ _11558_ keylen _10371_ _03341_ _03345_ sky130_fd_sc_hd__o221ai_2
X_11668_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[1\] dec_new_block\[1\]
+ _07398_ sky130_fd_sc_hd__mux2_2
XFILLER_0_86_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_944 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_98_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13407_ VGND VPWR VGND VPWR _08886_ _07712_ keymem.key_mem\[6\]\[124\] _08885_ _08020_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_52_752 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17175_ VPWR VGND VPWR VGND _03284_ key[75] _11109_ sky130_fd_sc_hd__or2_2
XFILLER_0_261_1108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14387_ VPWR VGND VPWR VGND _09854_ _09856_ _09857_ _09516_ _09853_ sky130_fd_sc_hd__or4b_2
XFILLER_0_113_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16126_ VGND VPWR VGND VPWR _11564_ _11390_ _11580_ _11484_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_40_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13338_ VPWR VGND VPWR VGND _08823_ keymem.key_mem\[3\]\[117\] _07844_ keymem.key_mem\[6\]\[117\]
+ _07771_ _08824_ sky130_fd_sc_hd__a221o_2
XFILLER_0_40_958 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16057_ VGND VPWR VGND VPWR _11466_ _11296_ _11512_ _11253_ sky130_fd_sc_hd__a21oi_2
X_13269_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[110\] _07622_ keymem.key_mem\[4\]\[110\]
+ _07637_ _08762_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_126_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15008_ VGND VPWR _10472_ _10439_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_249_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1338 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19816_ VGND VPWR VPWR VGND _05314_ keymem.key_mem\[11\]\[66\] _03209_ _05318_ sky130_fd_sc_hd__mux2_2
XFILLER_0_97_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19747_ VGND VPWR VPWR VGND _05281_ keymem.key_mem\[11\]\[33\] _02883_ _05282_ sky130_fd_sc_hd__mux2_2
X_16959_ VGND VPWR VGND VPWR _03089_ _03087_ _03086_ _09534_ _03088_ _09514_ sky130_fd_sc_hd__a32o_2
XFILLER_0_159_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_95_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19678_ VGND VPWR VPWR VGND _05243_ keymem.key_mem\[11\]\[1\] _09725_ _05245_ sky130_fd_sc_hd__mux2_2
XFILLER_0_220_920 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_204_Left_471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_154_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_133_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18629_ VPWR VGND _04497_ _04496_ enc_block.block_w1_reg\[28\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_137_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Right_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_231_290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_34_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21640_ VGND VPWR VPWR VGND _06286_ _02688_ keymem.key_mem\[4\]\[24\] _06288_ sky130_fd_sc_hd__mux2_2
XFILLER_0_136_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21571_ VGND VPWR VPWR VGND _06242_ _03627_ keymem.key_mem\[5\]\[121\] _06250_ sky130_fd_sc_hd__mux2_2
XFILLER_0_69_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23310_ VPWR VGND _07191_ _07190_ enc_block.round_key\[10\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_20522_ VGND VPWR VPWR VGND _05692_ _11039_ keymem.key_mem\[8\]\[13\] _05693_ sky130_fd_sc_hd__mux2_2
XFILLER_0_248_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24290_ VGND VPWR VPWR VGND clk _00783_ reset_n keymem.key_mem\[10\]\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_170_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_69_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23241_ VPWR VGND _07128_ enc_block.block_w2_reg\[7\] enc_block.block_w2_reg\[3\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_248_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20453_ VGND VPWR _00993_ _05655_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_213_Left_480 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23172_ VGND VPWR _02296_ _07071_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20384_ VGND VPWR _00960_ _05619_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_109_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22123_ VGND VPWR VPWR VGND _06538_ _05079_ keymem.key_mem\[3\]\[122\] _06545_ sky130_fd_sc_hd__mux2_2
XFILLER_0_112_161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1074 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_100_334 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_208_Right_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22054_ VGND VPWR VPWR VGND _06494_ _05015_ keymem.key_mem\[3\]\[89\] _06509_ sky130_fd_sc_hd__mux2_2
XFILLER_0_246_338 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_105_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21005_ VGND VPWR _01250_ _05950_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_103_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25813_ VGND VPWR VPWR VGND clk _02306_ reset_n enc_block.block_w3_reg\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_242_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_255_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25744_ keymem.prev_key1_reg\[60\] clk _02237_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22956_ VGND VPWR VGND VPWR _06941_ _02888_ _03860_ _06884_ _02892_ sky130_fd_sc_hd__a211o_2
XFILLER_0_186_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21907_ VGND VPWR VGND VPWR _06430_ keymem.key_mem_we _02480_ _06420_ _01672_ sky130_fd_sc_hd__a31o_2
XFILLER_0_214_1132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25675_ VGND VPWR VPWR VGND clk _02168_ reset_n keymem.rcon_logic.tmp_rcon\[5\] sky130_fd_sc_hd__dfrtp_2
X_22887_ VGND VPWR _10660_ keylen _06898_ _10382_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_116_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12640_ VPWR VGND VPWR VGND _08194_ keymem.key_mem\[5\]\[48\] _07811_ keymem.key_mem\[11\]\[48\]
+ _07781_ _08195_ sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_217_Right_86 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24626_ VGND VPWR VPWR VGND clk _01119_ reset_n keymem.key_mem\[8\]\[107\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_52_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21838_ VGND VPWR _01642_ _06391_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_210_1007 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_194_153 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_194_175 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_186_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12571_ VPWR VGND VPWR VGND _08132_ keymem.key_mem\[14\]\[41\] _07666_ keymem.key_mem\[2\]\[41\]
+ _08131_ _08133_ sky130_fd_sc_hd__a221o_2
X_24557_ VGND VPWR VPWR VGND clk _01050_ reset_n keymem.key_mem\[8\]\[38\] sky130_fd_sc_hd__dfrtp_2
X_21769_ VGND VPWR _06355_ _06258_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14310_ VPWR VGND VGND VPWR _09489_ _09780_ _09426_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_359 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23508_ VPWR VGND VPWR VGND aes_core_ctrl_reg\[0\] reset_n _00004_ clk sky130_fd_sc_hd__dfstp_2
X_15290_ VPWR VGND VGND VPWR _10565_ _10520_ _10752_ _10618_ _10751_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_80_324 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_266_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24488_ VGND VPWR VPWR VGND clk _00981_ reset_n keymem.key_mem\[9\]\[97\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_260_Right_129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14241_ VGND VPWR _09712_ keymem.prev_key0_reg\[33\] keymem.prev_key0_reg\[65\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
X_23439_ VGND VPWR _07306_ enc_block.block_w2_reg\[0\] _07157_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_227_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_774 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14172_ VGND VPWR VGND VPWR _09210_ _09096_ _09085_ _09050_ _09643_ sky130_fd_sc_hd__o22a_2
XFILLER_0_81_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13123_ VGND VPWR VGND VPWR _08631_ _07968_ keymem.key_mem\[9\]\[95\] _08628_ _08630_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_238_806 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25109_ VGND VPWR VPWR VGND clk _01602_ reset_n keymem.key_mem\[4\]\[78\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_226_Right_95 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18980_ VPWR VGND _04813_ _04812_ enc_block.round_key\[55\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_103_183 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_123_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17931_ VGND VPWR VPWR VGND _03876_ key[229] keymem.prev_key1_reg\[101\] _03885_
+ sky130_fd_sc_hd__mux2_2
X_13054_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[89\] _07743_ keymem.key_mem\[8\]\[89\]
+ _08211_ _08568_ sky130_fd_sc_hd__a22o_2
X_12005_ VGND VPWR enc_block.round_key\[0\] _07607_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_203_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_246_861 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17862_ VGND VPWR VGND VPWR _03316_ keymem.prev_key1_reg\[79\] _03838_ _03818_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_218_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19601_ VGND VPWR VPWR VGND _05183_ _05021_ keymem.key_mem\[12\]\[94\] _05203_ sky130_fd_sc_hd__mux2_2
X_16813_ VGND VPWR _00052_ _02956_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17793_ VPWR VGND VGND VPWR _03790_ _03791_ _03731_ sky130_fd_sc_hd__nor2_2
X_19532_ VPWR VGND keymem.key_mem\[12\]\[61\] _05167_ _05158_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16744_ VGND VPWR _02894_ _02893_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13956_ VGND VPWR VPWR VGND _09416_ _09415_ _09428_ _09427_ _09424_ sky130_fd_sc_hd__o211a_2
XFILLER_0_261_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_152_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_202_931 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19463_ VPWR VGND keymem.key_mem\[12\]\[29\] _05130_ _05128_ VPWR VGND sky130_fd_sc_hd__and2_2
X_12907_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[74\] _07651_ keymem.key_mem\[12\]\[74\]
+ _07673_ _08436_ sky130_fd_sc_hd__a22o_2
X_13887_ VPWR VGND VGND VPWR _09350_ _09353_ _09359_ _09358_ _09355_ sky130_fd_sc_hd__o22ai_2
X_16675_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[126\] _02818_ _02829_ _02819_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_92_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_158_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18414_ VGND VPWR _04303_ enc_block.sword_ctr_reg\[0\] _00306_ _04073_ VPWR VGND
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_124_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15626_ VGND VPWR VGND VPWR _10521_ _10546_ _10510_ _10587_ _11084_ sky130_fd_sc_hd__o22a_2
XFILLER_0_29_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12838_ VPWR VGND VPWR VGND _08373_ keymem.key_mem\[14\]\[67\] _07583_ keymem.key_mem\[10\]\[67\]
+ _07561_ _08374_ sky130_fd_sc_hd__a221o_2
X_19394_ VGND VPWR _00499_ _05090_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_56_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18345_ VPWR VGND _04242_ _03960_ enc_block.block_w1_reg\[17\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_267_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15557_ VGND VPWR VPWR VGND _10525_ _10564_ _10450_ _11016_ sky130_fd_sc_hd__or3_2
XFILLER_0_56_354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12769_ VPWR VGND VPWR VGND _08311_ keymem.key_mem\[5\]\[60\] _08052_ keymem.key_mem\[9\]\[60\]
+ _07705_ _08312_ sky130_fd_sc_hd__a221o_2
XFILLER_0_51_1073 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_56_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_302 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14508_ VPWR VGND VGND VPWR _09168_ _09687_ _09146_ _09107_ _09977_ _09976_ sky130_fd_sc_hd__o221a_2
X_15488_ VGND VPWR VGND VPWR _10924_ _10948_ _10935_ _10947_ _10930_ sky130_fd_sc_hd__and4bb_2
X_18276_ VPWR VGND VGND VPWR _04179_ _04180_ _04041_ sky130_fd_sc_hd__nor2_2
XFILLER_0_126_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_176_1_Right_777 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_83_195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17227_ VGND VPWR VPWR VGND _03296_ keymem.key_mem\[14\]\[80\] _03330_ _03331_ sky130_fd_sc_hd__mux2_2
X_14439_ VGND VPWR VPWR VGND _09905_ _09368_ _09908_ _09907_ _09906_ sky130_fd_sc_hd__o211a_2
XFILLER_0_64_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1047 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17158_ VGND VPWR VPWR VGND _03185_ keymem.key_mem\[14\]\[73\] _03268_ _03269_ sky130_fd_sc_hd__mux2_2
XFILLER_0_163_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16109_ VGND VPWR VGND VPWR _11562_ _11563_ _11482_ _11241_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_12_468 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_60_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17089_ VPWR VGND VPWR VGND _03207_ key[66] _09987_ sky130_fd_sc_hd__or2_2
XFILLER_0_0_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_625 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_58_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_490 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_58_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_850 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_58_1205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_251_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_100_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22810_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[111\] _06858_ _06857_ _05056_ _02147_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_28_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_86 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23790_ VGND VPWR VPWR VGND clk _00283_ reset_n enc_block.block_w0_reg\[9\] sky130_fd_sc_hd__dfrtp_2
X_22741_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[65\] _06820_ _06819_ _04975_ _02101_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_174_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_181_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25460_ VGND VPWR VPWR VGND clk _01953_ reset_n keymem.key_mem\[1\]\[45\] sky130_fd_sc_hd__dfrtp_2
X_22672_ VGND VPWR _02060_ _06807_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_9_Left_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_176_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_59_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24411_ VGND VPWR VPWR VGND clk _00904_ reset_n keymem.key_mem\[9\]\[20\] sky130_fd_sc_hd__dfrtp_2
X_21623_ VGND VPWR VPWR VGND _06275_ _11446_ keymem.key_mem\[4\]\[16\] _06279_ sky130_fd_sc_hd__mux2_2
X_25391_ VGND VPWR VPWR VGND clk _01884_ reset_n keymem.key_mem\[2\]\[104\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_176_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_48_899 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_69_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_162 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24342_ VGND VPWR VPWR VGND clk _00835_ reset_n keymem.key_mem\[10\]\[79\] sky130_fd_sc_hd__dfrtp_2
X_21554_ VGND VPWR VPWR VGND _06231_ _03573_ keymem.key_mem\[5\]\[113\] _06241_ sky130_fd_sc_hd__mux2_2
XFILLER_0_248_1250 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_209_1201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_191_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20505_ VGND VPWR VPWR VGND _05680_ _10193_ keymem.key_mem\[8\]\[5\] _05684_ sky130_fd_sc_hd__mux2_2
X_24273_ VGND VPWR VPWR VGND clk _00766_ reset_n keymem.key_mem\[10\]\[10\] sky130_fd_sc_hd__dfrtp_2
X_21485_ VGND VPWR VPWR VGND _06196_ _03329_ keymem.key_mem\[5\]\[80\] _06205_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_774 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23224_ VGND VPWR _07113_ enc_block.round_key\[2\] _07112_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20436_ VGND VPWR _00985_ _05646_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_209_1289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_181_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_766 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23155_ VGND VPWR VGND VPWR _07062_ _03562_ _06890_ _06924_ _03566_ sky130_fd_sc_hd__a211o_2
X_20367_ VGND VPWR _05610_ _03227_ _00952_ _05532_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_259_474 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22106_ VGND VPWR VPWR VGND _06527_ _05062_ keymem.key_mem\[3\]\[114\] _06536_ sky130_fd_sc_hd__mux2_2
XFILLER_0_179_1311 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23086_ VGND VPWR VGND VPWR _02263_ _07018_ _07010_ keymem.prev_key1_reg\[86\] sky130_fd_sc_hd__o21a_2
XFILLER_0_140_1145 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20298_ VGND VPWR _00919_ _05574_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22037_ VGND VPWR VGND VPWR _06500_ keymem.key_mem_we _03330_ _06498_ _01732_ sky130_fd_sc_hd__a31o_2
XFILLER_0_179_1355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_100_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_209_79 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_216_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13810_ VGND VPWR VGND VPWR _09282_ enc_block.block_w2_reg\[29\] enc_block.sword_ctr_reg\[1\]
+ enc_block.sword_ctr_reg\[0\] sky130_fd_sc_hd__and3b_2
X_14790_ VPWR VGND VPWR VGND _09247_ _09390_ _09425_ _09361_ _10256_ sky130_fd_sc_hd__or4_2
XFILLER_0_192_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23988_ VGND VPWR VPWR VGND clk _00481_ reset_n keymem.key_mem\[13\]\[109\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_97_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13741_ VGND VPWR VGND VPWR _09213_ _09207_ _09106_ _09208_ _09212_ sky130_fd_sc_hd__a211o_2
XFILLER_0_199_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25727_ keymem.prev_key1_reg\[43\] clk _02220_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22939_ VGND VPWR VGND VPWR _02754_ _06928_ _02763_ _06931_ sky130_fd_sc_hd__a21o_2
X_16460_ VGND VPWR VGND VPWR _11235_ _11399_ _11252_ _11497_ _02621_ sky130_fd_sc_hd__o22a_2
X_13672_ VPWR VGND VPWR VGND _08963_ _09064_ _09017_ _08957_ _09144_ sky130_fd_sc_hd__or4_2
X_25658_ VGND VPWR VPWR VGND clk _02151_ reset_n keymem.key_mem\[0\]\[115\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_167_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_304 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15411_ VPWR VGND VGND VPWR _10446_ _10872_ _10672_ _10475_ sky130_fd_sc_hd__nor3b_2
X_12623_ VGND VPWR VGND VPWR _08180_ _07725_ keymem.key_mem\[5\]\[46\] _08177_ _08179_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_2_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16391_ VPWR VGND VGND VPWR _02365_ _02376_ _02553_ sky130_fd_sc_hd__or2b_2
X_24609_ VGND VPWR VPWR VGND clk _01102_ reset_n keymem.key_mem\[8\]\[90\] sky130_fd_sc_hd__dfrtp_2
X_25589_ VGND VPWR VPWR VGND clk _02082_ reset_n keymem.key_mem\[0\]\[46\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_888 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15342_ VGND VPWR VGND VPWR _10562_ _10804_ _10464_ _10472_ _10459_ sky130_fd_sc_hd__and4bb_2
X_18130_ VGND VPWR _04046_ enc_block.block_w0_reg\[30\] _04045_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_87_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12554_ VPWR VGND VPWR VGND keymem.key_mem\[8\]\[40\] _07958_ keymem.key_mem\[2\]\[40\]
+ _08116_ _08117_ sky130_fd_sc_hd__a22o_2
XFILLER_0_54_858 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_1033 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_54_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_170_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18061_ VGND VPWR _03982_ _03981_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15273_ VGND VPWR VPWR VGND _10736_ _10731_ _10665_ _10735_ _09931_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_48_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12485_ VGND VPWR VGND VPWR _08055_ _08050_ keymem.key_mem\[7\]\[33\] _08051_ _08054_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_227_1345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_571 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14224_ VGND VPWR VGND VPWR _09145_ _09091_ _09695_ _09148_ sky130_fd_sc_hd__a21oi_2
X_17012_ VPWR VGND VPWR VGND _03137_ key[187] _10286_ sky130_fd_sc_hd__or2_2
XFILLER_0_21_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14155_ VPWR VGND VGND VPWR _09495_ _09422_ _09626_ _09311_ _09418_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_22_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1006 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13106_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[94\] _07782_ keymem.key_mem\[2\]\[94\]
+ _08116_ _08615_ sky130_fd_sc_hd__a22o_2
X_14086_ VPWR VGND VPWR VGND _09554_ _09556_ _09555_ _09551_ _09557_ sky130_fd_sc_hd__or4_2
X_18963_ VPWR VGND VPWR VGND _04797_ _04788_ _04796_ enc_block.block_w2_reg\[21\]
+ _04709_ _00361_ sky130_fd_sc_hd__a221o_2
XFILLER_0_197_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17914_ VGND VPWR VPWR VGND _03812_ key[224] keymem.prev_key1_reg\[96\] _03873_ sky130_fd_sc_hd__mux2_2
XFILLER_0_253_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13037_ VGND VPWR VGND VPWR _07808_ keymem.key_mem\[12\]\[87\] _08550_ _08552_ _08553_
+ _08480_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_266_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18894_ VGND VPWR VGND VPWR _04734_ _03992_ _04735_ _00354_ sky130_fd_sc_hd__a21o_2
XFILLER_0_98_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17845_ VGND VPWR _00214_ _03826_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_238_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17776_ VGND VPWR _00192_ _03779_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14988_ VGND VPWR VGND VPWR _10452_ _10401_ _10400_ keymem.prev_key1_reg\[10\] _08954_
+ _08941_ sky130_fd_sc_hd__a32o_2
XFILLER_0_261_694 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19515_ VGND VPWR VGND VPWR _05157_ keymem.key_mem_we _03083_ _05135_ _00553_ sky130_fd_sc_hd__a31o_2
X_16727_ VGND VPWR VGND VPWR _02878_ _10328_ _02877_ key[33] sky130_fd_sc_hd__o21a_2
XFILLER_0_260_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13939_ VGND VPWR _09411_ _09410_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_44_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1040 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19446_ VGND VPWR VGND VPWR _05120_ keymem.key_mem_we _02550_ _05109_ _00521_ sky130_fd_sc_hd__a31o_2
X_16658_ VGND VPWR VPWR VGND _02662_ keymem.key_mem\[14\]\[29\] _02812_ _02813_ sky130_fd_sc_hd__mux2_2
X_15609_ VGND VPWR VGND VPWR _10489_ _10513_ _10595_ _10583_ _11067_ sky130_fd_sc_hd__o22a_2
XFILLER_0_9_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_102_1_Left_369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19377_ VPWR VGND keymem.key_mem_we _05079_ _03633_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_17_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16589_ VGND VPWR VGND VPWR _02393_ _02372_ _02745_ _02746_ sky130_fd_sc_hd__a21o_2
XFILLER_0_151_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_169_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_527 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18328_ VGND VPWR _04227_ enc_block.block_w2_reg\[14\] enc_block.block_w2_reg\[15\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18259_ VPWR VGND VPWR VGND _04164_ _04162_ _04163_ sky130_fd_sc_hd__or2_2
XFILLER_0_154_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_177_1_Right_778 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_71_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_206_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21270_ VGND VPWR VPWR VGND _06087_ _03538_ keymem.key_mem\[6\]\[107\] _06091_ sky130_fd_sc_hd__mux2_2
XFILLER_0_206_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_1204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20221_ VPWR VGND VPWR VGND _05533_ _05532_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_164_1_Left_431 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_100_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_12_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_2_Left_603 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Right_4 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_106_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20152_ VGND VPWR VPWR VGND _05493_ _03466_ keymem.key_mem\[10\]\[96\] _05496_ sky130_fd_sc_hd__mux2_2
XFILLER_0_176_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24960_ VGND VPWR VPWR VGND clk _01453_ reset_n keymem.key_mem\[5\]\[57\] sky130_fd_sc_hd__dfrtp_2
X_20083_ VGND VPWR VPWR VGND _05457_ _03184_ keymem.key_mem\[10\]\[63\] _05460_ sky130_fd_sc_hd__mux2_2
XFILLER_0_228_179 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23911_ VGND VPWR VPWR VGND clk _00404_ reset_n keymem.key_mem\[13\]\[32\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_209_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_256_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24891_ VGND VPWR VPWR VGND clk _01384_ reset_n keymem.key_mem\[6\]\[116\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_252_661 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23842_ VGND VPWR VPWR VGND clk _00335_ reset_n enc_block.block_w1_reg\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_217_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23773_ VGND VPWR VPWR VGND clk _00008_ reset_n enc_block.sword_ctr_inc sky130_fd_sc_hd__dfrtp_2
XFILLER_0_135_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20985_ VGND VPWR VPWR VGND _05934_ _05035_ keymem.key_mem\[7\]\[101\] _05940_ sky130_fd_sc_hd__mux2_2
XFILLER_0_71_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_192_95 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22724_ VGND VPWR VPWR VGND _06822_ keymem.key_mem\[0\]\[57\] _03119_ _06827_ sky130_fd_sc_hd__mux2_2
X_25512_ VGND VPWR VPWR VGND clk _02005_ reset_n keymem.key_mem\[1\]\[97\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_152_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_71_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1184 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25443_ VGND VPWR VPWR VGND clk _01936_ reset_n keymem.key_mem\[1\]\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_137_315 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_36_803 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22655_ VGND VPWR VPWR VGND _06798_ keymem.key_mem\[0\]\[16\] _11447_ _06799_ sky130_fd_sc_hd__mux2_2
XFILLER_0_137_326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_164_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_47_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21606_ VGND VPWR VPWR VGND _06263_ _10661_ keymem.key_mem\[4\]\[8\] _06270_ sky130_fd_sc_hd__mux2_2
X_25374_ VGND VPWR VPWR VGND clk _01867_ reset_n keymem.key_mem\[2\]\[87\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_8_760 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22586_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[100\] _06767_ _06766_ _05033_ _02008_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_36_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_127_2_Left_598 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_111_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24325_ VGND VPWR VPWR VGND clk _00818_ reset_n keymem.key_mem\[10\]\[62\] sky130_fd_sc_hd__dfrtp_2
X_21537_ VGND VPWR _01500_ _06232_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_62_176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_96_1_Left_363 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12270_ VGND VPWR VGND VPWR _07858_ _07731_ keymem.key_mem\[13\]\[15\] _07853_ _07857_
+ sky130_fd_sc_hd__a211o_2
X_24256_ VGND VPWR VPWR VGND clk _00749_ reset_n keymem.key_mem\[11\]\[121\] sky130_fd_sc_hd__dfrtp_2
X_21468_ VGND VPWR _06196_ _06115_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_82_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23207_ VGND VPWR _07097_ enc_block.block_w1_reg\[9\] _07086_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_146_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20419_ VGND VPWR _00977_ _05637_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_120_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24187_ VGND VPWR VPWR VGND clk _00680_ reset_n keymem.key_mem\[11\]\[52\] sky130_fd_sc_hd__dfrtp_2
X_21399_ VGND VPWR VPWR VGND _06151_ _02945_ keymem.key_mem\[5\]\[39\] _06160_ sky130_fd_sc_hd__mux2_2
XFILLER_0_31_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_82_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23138_ VGND VPWR VPWR VGND _07032_ _07050_ keymem.prev_key1_reg\[106\] _07051_ sky130_fd_sc_hd__mux2_2
XFILLER_0_208_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_189_2_Left_660 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15960_ VPWR VGND VGND VPWR _11270_ _11327_ _11416_ _11182_ _11330_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_41_1050 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23069_ VGND VPWR VPWR VGND _02256_ _03317_ _03320_ _06976_ _07008_ sky130_fd_sc_hd__o31a_2
XPHY_EDGE_ROW_139_1_Right_740 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14911_ VGND VPWR keymem.prev_key1_reg\[72\] _10373_ _10375_ _10374_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_15891_ VGND VPWR VGND VPWR _11303_ _11257_ _11347_ _11280_ sky130_fd_sc_hd__a21oi_2
X_17630_ VGND VPWR _00143_ _03682_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14842_ VGND VPWR VGND VPWR _09415_ _09302_ _09391_ _09478_ _09437_ _10307_ sky130_fd_sc_hd__o32a_2
XFILLER_0_76_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17561_ VGND VPWR VGND VPWR _02710_ _02709_ _03624_ _10967_ sky130_fd_sc_hd__a21oi_2
X_14773_ VGND VPWR VPWR VGND _09564_ _09392_ _10239_ _10238_ _09742_ sky130_fd_sc_hd__o211a_2
XFILLER_0_93_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11985_ VGND VPWR _07588_ _07587_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_153_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19300_ VPWR VGND keymem.key_mem_we _05027_ _03474_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16512_ VPWR VGND VGND VPWR _02672_ _02667_ _02671_ sky130_fd_sc_hd__nand2_2
X_13724_ VPWR VGND VGND VPWR _09196_ _09041_ _09040_ sky130_fd_sc_hd__nand2_2
X_17492_ VPWR VGND VGND VPWR _03564_ key[240] _10278_ sky130_fd_sc_hd__nand2_2
XFILLER_0_54_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_39_641 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_252_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19231_ VGND VPWR _00442_ _04984_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16443_ VGND VPWR VGND VPWR _02603_ _02601_ _02605_ _02604_ sky130_fd_sc_hd__a21oi_2
X_13655_ VGND VPWR _09127_ _09126_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_195_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12606_ VGND VPWR enc_block.round_key\[44\] _08164_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19162_ VGND VPWR _00415_ _04942_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13586_ VGND VPWR _09058_ _09030_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16374_ VPWR VGND VPWR VGND _02536_ _02537_ _07385_ _02498_ sky130_fd_sc_hd__or3b_2
XFILLER_0_186_1145 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18113_ VGND VPWR VPWR VGND _03974_ enc_block.block_w0_reg\[4\] _04030_ _04031_ sky130_fd_sc_hd__mux2_2
X_15325_ VGND VPWR VGND VPWR _10509_ _10414_ _10787_ _10540_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_53_143 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12537_ VGND VPWR VGND VPWR _08102_ _07854_ keymem.key_mem\[4\]\[38\] _08101_ _07746_
+ sky130_fd_sc_hd__a211o_2
X_19093_ VPWR VGND keymem.key_mem\[13\]\[16\] _04901_ _04887_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_41_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18044_ VGND VPWR _03966_ _03965_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_164_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15256_ VPWR VGND VPWR VGND _10719_ _10562_ _10718_ sky130_fd_sc_hd__or2_2
X_12468_ VPWR VGND VPWR VGND _08038_ keymem.key_mem\[13\]\[32\] _07730_ keymem.key_mem\[14\]\[32\]
+ _07706_ _08039_ sky130_fd_sc_hd__a221o_2
XFILLER_0_2_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_160_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14207_ VPWR VGND VPWR VGND _09678_ _09198_ _09048_ sky130_fd_sc_hd__or2_2
XFILLER_0_164_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15187_ VPWR VGND VPWR VGND _10643_ _10650_ _10648_ _10637_ _10651_ sky130_fd_sc_hd__or4_2
X_12399_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[26\] _07564_ keymem.key_mem\[2\]\[26\]
+ _07545_ _07976_ sky130_fd_sc_hd__a22o_2
XFILLER_0_240_1331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14138_ VGND VPWR VGND VPWR _09437_ _09430_ _09318_ _09410_ _09609_ sky130_fd_sc_hd__o22a_2
XFILLER_0_61_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19995_ VGND VPWR VPWR VGND _05413_ _02550_ keymem.key_mem\[10\]\[21\] _05414_ sky130_fd_sc_hd__mux2_2
XFILLER_0_254_915 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_190_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18946_ VGND VPWR _04782_ enc_block.block_w1_reg\[4\] enc_block.block_w0_reg\[12\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_14069_ VGND VPWR _09541_ _09540_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_253_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18877_ VPWR VGND VPWR VGND _04720_ enc_block.block_w1_reg\[4\] enc_block.block_w1_reg\[5\]
+ sky130_fd_sc_hd__or2_2
XFILLER_0_101_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17828_ VGND VPWR VPWR VGND _03814_ _03813_ keymem.prev_key0_reg\[68\] _03815_ sky130_fd_sc_hd__mux2_2
XFILLER_0_171_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17759_ VGND VPWR VPWR VGND _03719_ key[172] keymem.prev_key1_reg\[44\] _03770_ sky130_fd_sc_hd__mux2_2
XFILLER_0_171_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1090 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_72_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20770_ VGND VPWR VGND VPWR _05825_ keymem.key_mem_we _09537_ _05821_ _01140_ sky130_fd_sc_hd__a31o_2
XFILLER_0_18_1085 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_251_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19429_ VGND VPWR VGND VPWR _05111_ keymem.key_mem_we _11040_ _05109_ _00513_ sky130_fd_sc_hd__a31o_2
XFILLER_0_91_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_212_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_186_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22440_ VGND VPWR _01922_ _06713_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_18_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_95_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22371_ VGND VPWR _01890_ _06676_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_44_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24110_ VGND VPWR VPWR VGND clk _00603_ reset_n keymem.key_mem\[12\]\[103\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_636 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21322_ VGND VPWR VPWR VGND _06117_ _09861_ keymem.key_mem\[5\]\[2\] _06120_ sky130_fd_sc_hd__mux2_2
X_25090_ VGND VPWR VPWR VGND clk _01583_ reset_n keymem.key_mem\[4\]\[59\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_182_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_349 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_178_1_Right_779 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24041_ VGND VPWR VPWR VGND clk _00534_ reset_n keymem.key_mem\[12\]\[34\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_143_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21253_ VGND VPWR VPWR VGND _06076_ _03485_ keymem.key_mem\[6\]\[99\] _06082_ sky130_fd_sc_hd__mux2_2
XFILLER_0_40_360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_1061 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_64_1083 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20204_ VGND VPWR VPWR VGND _05515_ _03627_ keymem.key_mem\[10\]\[121\] _05523_ sky130_fd_sc_hd__mux2_2
X_21184_ VGND VPWR VPWR VGND _06040_ _03209_ keymem.key_mem\[6\]\[66\] _06046_ sky130_fd_sc_hd__mux2_2
X_20135_ VGND VPWR VPWR VGND _05482_ _03401_ keymem.key_mem\[10\]\[88\] _05487_ sky130_fd_sc_hd__mux2_2
XFILLER_0_217_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_99_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_447 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20066_ VGND VPWR VPWR VGND _05446_ _03099_ keymem.key_mem\[10\]\[55\] _05451_ sky130_fd_sc_hd__mux2_2
XFILLER_0_239_1046 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24943_ VGND VPWR VPWR VGND clk _01436_ reset_n keymem.key_mem\[5\]\[40\] sky130_fd_sc_hd__dfrtp_2
X_24874_ VGND VPWR VPWR VGND clk _01367_ reset_n keymem.key_mem\[6\]\[99\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_213_834 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23825_ VGND VPWR VPWR VGND clk _00318_ reset_n enc_block.block_w1_reg\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_240_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_169_259 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_240_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11770_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[20\] dec_new_block\[52\]
+ _07449_ sky130_fd_sc_hd__mux2_2
X_23756_ keymem.prev_key0_reg\[112\] clk _00253_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20968_ VPWR VGND keymem.key_mem\[7\]\[93\] _05931_ _05823_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_230_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_67_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22707_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[46\] _06820_ _06819_ _04947_ _02082_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_215_1090 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23687_ keymem.prev_key0_reg\[43\] clk _00184_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20899_ VPWR VGND keymem.key_mem\[7\]\[60\] _05895_ _05886_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_230_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13440_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[127\] _07666_ keymem.key_mem\[10\]\[127\]
+ _07876_ _08916_ sky130_fd_sc_hd__a22o_2
XFILLER_0_82_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22638_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[7\] _06790_ _06789_ _04889_ _02043_
+ sky130_fd_sc_hd__a22o_2
X_25426_ VGND VPWR VPWR VGND clk _01919_ reset_n keymem.key_mem\[1\]\[11\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_36_633 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_64_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25357_ VGND VPWR VPWR VGND clk _01850_ reset_n keymem.key_mem\[2\]\[70\] sky130_fd_sc_hd__dfrtp_2
X_13371_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[120\] _08391_ keymem.key_mem\[14\]\[120\]
+ _07744_ _08854_ sky130_fd_sc_hd__a22o_2
X_22569_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[88\] _06767_ _06766_ _05013_ _01996_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_1_1172 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_50_102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1331 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15110_ VGND VPWR _10574_ _10573_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12322_ VGND VPWR VGND VPWR _07584_ keymem.key_mem\[14\]\[19\] _07898_ _07900_ _07906_
+ _07905_ sky130_fd_sc_hd__a2111o_2
X_16090_ VGND VPWR VPWR VGND _11542_ _11541_ _11545_ _09722_ _11544_ sky130_fd_sc_hd__o211a_2
X_24308_ VGND VPWR VPWR VGND clk _00801_ reset_n keymem.key_mem\[10\]\[45\] sky130_fd_sc_hd__dfrtp_2
X_25288_ VGND VPWR VPWR VGND clk _01781_ reset_n keymem.key_mem\[2\]\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_224_1326 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15041_ VGND VPWR VGND VPWR _10502_ _10501_ _10505_ _10504_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_133_384 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12253_ VGND VPWR _07842_ _07705_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24239_ VGND VPWR VPWR VGND clk _00732_ reset_n keymem.key_mem\[11\]\[104\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_239_219 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_47_1270 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12184_ VPWR VGND VPWR VGND _07776_ keymem.key_mem\[8\]\[10\] _07753_ keymem.key_mem\[2\]\[10\]
+ _07547_ _07777_ sky130_fd_sc_hd__a221o_2
XFILLER_0_236_904 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_222_1061 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18800_ _04649_ _04651_ _04560_ _04650_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_248_775 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_101_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19780_ VGND VPWR VPWR VGND _05292_ keymem.key_mem\[11\]\[49\] _03046_ _05299_ sky130_fd_sc_hd__mux2_2
XFILLER_0_263_723 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16992_ VGND VPWR _03119_ _03118_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_78_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18731_ VPWR VGND VPWR VGND _04587_ block[95] _04576_ enc_block.block_w1_reg\[31\]
+ _04543_ _04588_ sky130_fd_sc_hd__a221o_2
X_15943_ VGND VPWR _11399_ _11398_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_250_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18662_ VPWR VGND _04527_ _04526_ enc_block.round_key\[87\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_92_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15874_ VGND VPWR _11330_ _11329_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17613_ VGND VPWR _00139_ _03669_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14825_ VGND VPWR VGND VPWR _10290_ _09785_ _09782_ _09560_ _09558_ sky130_fd_sc_hd__and4_2
XFILLER_0_157_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18593_ _04463_ _04465_ _04064_ _04464_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_98_360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_230_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_204_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17544_ VGND VPWR VPWR VGND _03029_ _03388_ key[119] _03609_ sky130_fd_sc_hd__mux2_2
X_14756_ VPWR VGND VPWR VGND _10217_ _10221_ _10222_ _10178_ _10181_ sky130_fd_sc_hd__or4b_2
X_11968_ VPWR VGND VGND VPWR _07527_ _07530_ _07571_ _07532_ _07531_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_15_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_153_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13707_ VPWR VGND VGND VPWR _09178_ _09179_ _09177_ sky130_fd_sc_hd__nor2_2
X_17475_ VPWR VGND VPWR VGND _03549_ _03494_ _03546_ key[237] _03527_ _03550_ sky130_fd_sc_hd__a221o_2
XFILLER_0_6_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14687_ VPWR VGND VGND VPWR _09114_ _10154_ _09687_ sky130_fd_sc_hd__nor2_2
XFILLER_0_73_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11899_ VGND VPWR result[116] _07513_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_132_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_15_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19214_ VPWR VGND keymem.key_mem\[13\]\[64\] _04974_ _04961_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16426_ VGND VPWR VGND VPWR _02588_ _02587_ _02552_ keymem.prev_key0_reg\[118\] sky130_fd_sc_hd__and3b_2
X_13638_ VGND VPWR _09110_ _09081_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_73_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19145_ VPWR VGND keymem.key_mem_we _04931_ _02934_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16357_ VGND VPWR VGND VPWR _11325_ _11527_ _11375_ _11385_ _02520_ sky130_fd_sc_hd__o22a_2
XFILLER_0_41_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13569_ VGND VPWR _09041_ _08970_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_203_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15308_ VGND VPWR VGND VPWR _10639_ _10541_ _10770_ _10769_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_41_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19076_ VGND VPWR VGND VPWR _04891_ keymem.key_mem_we _10662_ _04878_ _00380_ sky130_fd_sc_hd__a31o_2
X_16288_ VGND VPWR VGND VPWR _02452_ _11291_ _11432_ _11426_ _11348_ _11377_ sky130_fd_sc_hd__a32o_2
XFILLER_0_42_658 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_164_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_722 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_124_384 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18027_ VGND VPWR _03949_ _03948_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15239_ VPWR VGND VGND VPWR _10602_ _10702_ _10588_ sky130_fd_sc_hd__nor2_2
XFILLER_0_258_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_125_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_239_720 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_164_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_254 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_788 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_572 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1369 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_61_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19978_ VGND VPWR VPWR VGND _05400_ _11040_ keymem.key_mem\[10\]\[13\] _05405_ sky130_fd_sc_hd__mux2_2
XFILLER_0_66_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18929_ VPWR VGND VPWR VGND _04766_ block[50] _04744_ enc_block.block_w3_reg\[18\]
+ _04666_ _04767_ sky130_fd_sc_hd__a221o_2
XFILLER_0_254_778 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_235_970 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21940_ VGND VPWR VGND VPWR _06448_ keymem.key_mem_we _02904_ _06446_ _01687_ sky130_fd_sc_hd__a31o_2
XFILLER_0_173_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_136_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21871_ VPWR VGND keymem.key_mem\[3\]\[4\] _06411_ _06406_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_175_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23610_ VGND VPWR VPWR VGND clk _00111_ reset_n keymem.key_mem\[14\]\[99\] sky130_fd_sc_hd__dfrtp_2
X_20822_ VGND VPWR VGND VPWR _05853_ keymem.key_mem_we _02689_ _05850_ _01164_ sky130_fd_sc_hd__a31o_2
XFILLER_0_171_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24590_ VGND VPWR VPWR VGND clk _01083_ reset_n keymem.key_mem\[8\]\[71\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_72_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23541_ VGND VPWR VPWR VGND clk _00042_ reset_n keymem.key_mem\[14\]\[30\] sky130_fd_sc_hd__dfrtp_2
X_20753_ VGND VPWR _01135_ _05813_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_159_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_33_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23472_ VPWR VGND _07335_ enc_block.block_w0_reg\[20\] enc_block.block_w2_reg\[4\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_20684_ VGND VPWR _01102_ _05777_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_134_104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25211_ VGND VPWR VPWR VGND clk _01704_ reset_n keymem.key_mem\[3\]\[52\] sky130_fd_sc_hd__dfrtp_2
X_22423_ VGND VPWR VPWR VGND _06702_ keymem.key_mem\[1\]\[6\] _10284_ _06705_ sky130_fd_sc_hd__mux2_2
X_25142_ VGND VPWR VPWR VGND clk _01635_ reset_n keymem.key_mem\[4\]\[111\] sky130_fd_sc_hd__dfrtp_2
X_22354_ VGND VPWR _01882_ _06667_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_66_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_147_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_861 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21305_ VGND VPWR VPWR VGND _05971_ _03647_ keymem.key_mem\[6\]\[124\] _06109_ sky130_fd_sc_hd__mux2_2
XFILLER_0_60_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25073_ VGND VPWR VPWR VGND clk _01566_ reset_n keymem.key_mem\[4\]\[42\] sky130_fd_sc_hd__dfrtp_2
X_22285_ VGND VPWR _01849_ _06631_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_44_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_143_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_680 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_182_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24024_ VGND VPWR VPWR VGND clk _00517_ reset_n keymem.key_mem\[12\]\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_104_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21236_ VGND VPWR VPWR VGND _06065_ _03426_ keymem.key_mem\[6\]\[91\] _06073_ sky130_fd_sc_hd__mux2_2
XFILLER_0_143_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_223_1370 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_257_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_40_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21167_ VGND VPWR VPWR VGND _06029_ _03129_ keymem.key_mem\[6\]\[58\] _06037_ sky130_fd_sc_hd__mux2_2
X_20118_ VGND VPWR VPWR VGND _05469_ _03330_ keymem.key_mem\[10\]\[80\] _05478_ sky130_fd_sc_hd__mux2_2
X_21098_ VGND VPWR VPWR VGND _05996_ _02720_ keymem.key_mem\[6\]\[25\] _06001_ sky130_fd_sc_hd__mux2_2
XFILLER_0_258_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_260_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20049_ VGND VPWR VPWR VGND _05435_ _03025_ keymem.key_mem\[10\]\[47\] _05442_ sky130_fd_sc_hd__mux2_2
X_12940_ VGND VPWR VGND VPWR _08466_ _08150_ keymem.key_mem\[3\]\[77\] _08463_ _08465_
+ sky130_fd_sc_hd__a211o_2
X_24926_ VGND VPWR VPWR VGND clk _01419_ reset_n keymem.key_mem\[5\]\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_244_299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_99_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_154_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12871_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[70\] _08259_ _08403_ _08399_ _08404_
+ sky130_fd_sc_hd__o22a_2
X_24857_ VGND VPWR VPWR VGND clk _01350_ reset_n keymem.key_mem\[6\]\[82\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_193_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_450 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_115_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_213_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_201_815 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14610_ VGND VPWR VGND VPWR _10076_ keymem.prev_key0_reg\[100\] _10078_ _10032_ sky130_fd_sc_hd__nand3_2
X_11822_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[14\] dec_new_block\[78\]
+ _07475_ sky130_fd_sc_hd__mux2_2
X_23808_ VGND VPWR VPWR VGND clk _00301_ reset_n enc_block.block_w0_reg\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_197_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15590_ VGND VPWR _11048_ _11044_ _11047_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24788_ VGND VPWR VPWR VGND clk _01281_ reset_n keymem.key_mem\[6\]\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_90_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11753_ VGND VPWR result[43] _07440_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14541_ VGND VPWR VGND VPWR _09012_ _09196_ _09705_ _10008_ _10009_ _09672_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_189_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_363 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23739_ keymem.prev_key0_reg\[95\] clk _00236_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_7_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17260_ VPWR VGND VPWR VGND _03360_ key[84] _08936_ sky130_fd_sc_hd__or2_2
XFILLER_0_113_1172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14472_ VPWR VGND VGND VPWR _09227_ _09669_ _09940_ _09941_ sky130_fd_sc_hd__nor3_2
X_11684_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[9\] dec_new_block\[9\]
+ _07406_ sky130_fd_sc_hd__mux2_2
X_16211_ VGND VPWR VGND VPWR _11283_ _11318_ _11404_ _11466_ _02376_ sky130_fd_sc_hd__o22a_2
XFILLER_0_265_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25409_ VGND VPWR VPWR VGND clk _01902_ reset_n keymem.key_mem\[2\]\[122\] sky130_fd_sc_hd__dfrtp_2
X_13423_ VGND VPWR VGND VPWR _08901_ _07665_ keymem.key_mem\[4\]\[125\] _08898_ _08900_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_3_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17191_ VPWR VGND VPWR VGND _03298_ keymem.prev_key0_reg\[77\] sky130_fd_sc_hd__inv_2
XFILLER_0_187_1295 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16142_ VPWR VGND VGND VPWR _11422_ _11596_ _11395_ sky130_fd_sc_hd__nor2_2
XFILLER_0_23_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13354_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[118\] _08027_ _08838_ _08832_ _08839_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_180_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12305_ VPWR VGND VPWR VGND _07889_ keymem.key_mem\[3\]\[18\] _07603_ keymem.key_mem\[6\]\[18\]
+ _07759_ _07890_ sky130_fd_sc_hd__a221o_2
XFILLER_0_165_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16073_ VGND VPWR VGND VPWR _11527_ _11239_ _11528_ _11460_ sky130_fd_sc_hd__a21oi_2
X_13285_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[111\] _07793_ _08776_ _08772_ enc_block.round_key\[111\]
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_133_192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_820 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15024_ VPWR VGND VPWR VGND _10473_ _10466_ _10453_ _10439_ _10488_ sky130_fd_sc_hd__or4_2
X_19901_ VGND VPWR _00734_ _05362_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12236_ VGND VPWR VGND VPWR _07799_ keymem.key_mem\[1\]\[13\] _07823_ _07825_ _07826_
+ _07572_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_122_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_258_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_387 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_241_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_915 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_259_Left_526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19832_ VPWR VGND VGND VPWR _05326_ keymem.key_mem\[11\]\[74\] _05243_ sky130_fd_sc_hd__nand2_2
XFILLER_0_196_1509 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12167_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[8\] _07596_ keymem.key_mem\[11\]\[8\]
+ _07761_ _07762_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_583 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_258_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_520 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_202_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_1_Left_378 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19763_ VGND VPWR VPWR VGND _05281_ keymem.key_mem\[11\]\[41\] _02964_ _05290_ sky130_fd_sc_hd__mux2_2
XFILLER_0_224_907 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12098_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[5\] _07695_ keymem.key_mem\[4\]\[5\]
+ _07693_ _07696_ sky130_fd_sc_hd__a22o_2
X_16975_ VGND VPWR VPWR VGND _03101_ _02691_ _03103_ _09514_ _03102_ sky130_fd_sc_hd__o211a_2
XFILLER_0_208_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_194_1244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18714_ VPWR VGND VPWR VGND _04572_ block[93] _04487_ enc_block.block_w1_reg\[29\]
+ _04543_ _04573_ sky130_fd_sc_hd__a221o_2
X_15926_ VGND VPWR VGND VPWR _11382_ _11378_ _11375_ _11311_ _11381_ sky130_fd_sc_hd__o211ai_2
X_19694_ VGND VPWR VPWR VGND _05247_ keymem.key_mem\[11\]\[8\] _10662_ _05254_ sky130_fd_sc_hd__mux2_2
XFILLER_0_36_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18645_ VGND VPWR _04512_ _04314_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15857_ VGND VPWR _11313_ _11312_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_172_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14808_ _10243_ _10274_ keymem.prev_key1_reg\[102\] _10261_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_188_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18576_ VPWR VGND _04450_ _04449_ enc_block.round_key\[78\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_172_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15788_ VPWR VGND VPWR VGND _11172_ _11216_ _11243_ _11232_ _11244_ sky130_fd_sc_hd__or4_2
XFILLER_0_133_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_173_1_Left_440 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17527_ VGND VPWR _00128_ _03594_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_15_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14739_ VGND VPWR VGND VPWR _09658_ _09222_ _09116_ _09157_ _10205_ sky130_fd_sc_hd__o22a_2
XFILLER_0_213_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_588 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_141_2_Left_612 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_200_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17458_ VGND VPWR _00118_ _03535_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_46_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_89_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16409_ VPWR VGND VGND VPWR _02571_ _02568_ _02570_ sky130_fd_sc_hd__nand2_2
XFILLER_0_116_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17389_ VGND VPWR _00109_ _03475_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_171_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_794 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19128_ VPWR VGND keymem.key_mem_we _04920_ _02873_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_131_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_171_298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_112_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19059_ VPWR VGND keymem.key_mem\[13\]\[1\] _04882_ _04880_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_124_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22070_ VGND VPWR _01748_ _06517_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_11_853 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_140_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21021_ VGND VPWR VPWR VGND _05956_ _05071_ keymem.key_mem\[7\]\[118\] _05959_ sky130_fd_sc_hd__mux2_2
XFILLER_0_11_886 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_58_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_881 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_239_572 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_542 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_242_726 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22972_ VGND VPWR VGND VPWR _06888_ keymem.prev_key1_reg\[40\] _06950_ _02217_ sky130_fd_sc_hd__o21ba_2
X_25760_ keymem.prev_key1_reg\[76\] clk _02253_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_78_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_184_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24711_ VGND VPWR VPWR VGND clk _01204_ reset_n keymem.key_mem\[7\]\[64\] sky130_fd_sc_hd__dfrtp_2
X_21923_ VGND VPWR _06439_ _06405_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25691_ keymem.prev_key1_reg\[7\] clk _02184_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_179_354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24642_ VGND VPWR VPWR VGND clk _01135_ reset_n keymem.key_mem\[8\]\[123\] sky130_fd_sc_hd__dfrtp_2
X_21854_ VGND VPWR _01650_ _06399_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_136_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_2_Left_544 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20805_ VGND VPWR _05844_ _05823_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_72_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21785_ VGND VPWR _01617_ _06363_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24573_ VGND VPWR VPWR VGND clk _01066_ reset_n keymem.key_mem\[8\]\[54\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_942 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20736_ VGND VPWR _01127_ _05804_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23524_ VGND VPWR VPWR VGND clk _00025_ reset_n keymem.key_mem\[14\]\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1093 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_92_355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23455_ VPWR VGND VPWR VGND _07320_ enc_block.block_w3_reg\[25\] enc_block.block_w1_reg\[10\]
+ sky130_fd_sc_hd__or2_2
X_20667_ VGND VPWR _01094_ _05768_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22406_ VGND VPWR _01907_ _06694_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23386_ VPWR VGND VPWR VGND _07259_ _07184_ _07257_ sky130_fd_sc_hd__or2_2
XFILLER_0_208_1129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_33_444 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_122_118 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20598_ VGND VPWR _01061_ _05732_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_225_1410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22337_ VGND VPWR VPWR VGND _06658_ _03452_ keymem.key_mem\[2\]\[94\] _06659_ sky130_fd_sc_hd__mux2_2
X_25125_ VGND VPWR VPWR VGND clk _01618_ reset_n keymem.key_mem\[4\]\[94\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_260_1334 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_60_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_347 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13070_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[90\] _08391_ keymem.key_mem\[9\]\[90\]
+ _07612_ _08583_ sky130_fd_sc_hd__a22o_2
X_25056_ VGND VPWR VPWR VGND clk _01549_ reset_n keymem.key_mem\[4\]\[25\] sky130_fd_sc_hd__dfrtp_2
X_22268_ VGND VPWR VPWR VGND _06622_ _03161_ keymem.key_mem\[2\]\[61\] _06623_ sky130_fd_sc_hd__mux2_2
XFILLER_0_237_509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24007_ VGND VPWR VPWR VGND clk _00500_ reset_n keymem.key_mem\[12\]\[0\] sky130_fd_sc_hd__dfrtp_2
X_12021_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[1\] _07622_ keymem.key_mem\[12\]\[1\]
+ _07621_ _07623_ sky130_fd_sc_hd__a22o_2
XFILLER_0_44_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21219_ VGND VPWR VPWR VGND _06052_ _03355_ keymem.key_mem\[6\]\[83\] _06064_ sky130_fd_sc_hd__mux2_2
X_22199_ VGND VPWR _01808_ _06586_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_79_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_512 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_233_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16760_ VGND VPWR _08927_ keymem.prev_key1_reg\[36\] _02908_ keymem.prev_key1_reg\[68\]
+ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_13972_ VGND VPWR _09444_ _09443_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15711_ VGND VPWR _11167_ _11166_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_232_247 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12923_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[76\] _07695_ keymem.key_mem\[1\]\[76\]
+ _07901_ _08450_ sky130_fd_sc_hd__a22o_2
X_24909_ VGND VPWR VPWR VGND clk _01402_ reset_n keymem.key_mem\[5\]\[6\] sky130_fd_sc_hd__dfrtp_2
X_16691_ VGND VPWR VPWR VGND _02841_ _02842_ keymem.rcon_logic.tmp_rcon\[0\] _02844_
+ sky130_fd_sc_hd__or3_2
X_18430_ VGND VPWR _04317_ _04316_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15642_ VGND VPWR VPWR VGND _11041_ keymem.key_mem\[14\]\[14\] _11099_ _11100_ sky130_fd_sc_hd__mux2_2
XFILLER_0_115_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12854_ VPWR VGND VPWR VGND _08387_ keymem.key_mem\[6\]\[69\] _07739_ keymem.key_mem\[10\]\[69\]
+ _07865_ _08388_ sky130_fd_sc_hd__a221o_2
XFILLER_0_154_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_706 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_197_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11805_ VGND VPWR result[69] _07466_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18361_ VPWR VGND VGND VPWR _04256_ _04257_ _04190_ sky130_fd_sc_hd__nor2_2
X_15573_ VGND VPWR keymem.prev_key1_reg\[77\] _11030_ _11032_ _11031_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_115_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12785_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[62\] _08125_ keymem.key_mem\[1\]\[62\]
+ _07671_ _08326_ sky130_fd_sc_hd__a22o_2
XFILLER_0_201_678 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_113_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17312_ VPWR VGND VGND VPWR _09732_ _03407_ key[217] sky130_fd_sc_hd__nor2_2
XFILLER_0_12_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14524_ VGND VPWR VPWR VGND _09864_ keymem.key_mem\[14\]\[3\] _09992_ _09993_ sky130_fd_sc_hd__mux2_2
X_18292_ VGND VPWR _04194_ _04118_ _04193_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11736_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[3\] dec_new_block\[35\]
+ _07432_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_344 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_138_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17243_ VPWR VGND VPWR VGND _03344_ _03345_ _10190_ _03343_ sky130_fd_sc_hd__or3b_2
XFILLER_0_153_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14455_ VPWR VGND VGND VPWR _09924_ _09883_ _09923_ sky130_fd_sc_hd__nand2_2
X_11667_ VGND VPWR result[0] _07397_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13406_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[124\] _08090_ keymem.key_mem\[10\]\[124\]
+ _07743_ _08885_ sky130_fd_sc_hd__a22o_2
X_17174_ VGND VPWR _03283_ keymem.prev_key0_reg\[75\] _03282_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_1140 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14386_ VGND VPWR _09856_ keymem.prev_key0_reg\[2\] _09855_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_226_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16125_ _11377_ _11579_ _11266_ _11357_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_3_349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_24_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13337_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[117\] _07631_ keymem.key_mem\[2\]\[117\]
+ _07545_ _08823_ sky130_fd_sc_hd__a22o_2
XFILLER_0_11_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_126_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16056_ VGND VPWR VPWR VGND _11507_ _11510_ _11505_ _11511_ sky130_fd_sc_hd__or3_2
XFILLER_0_121_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13268_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[110\] _07778_ keymem.key_mem\[6\]\[110\]
+ _07908_ _08761_ sky130_fd_sc_hd__a22o_2
XFILLER_0_122_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15007_ VPWR VGND VPWR VGND _10460_ _10470_ _10471_ _10438_ _10450_ sky130_fd_sc_hd__or4b_2
XFILLER_0_23_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12219_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[12\] _07652_ keymem.key_mem\[11\]\[12\]
+ _07809_ _07810_ sky130_fd_sc_hd__a22o_2
XFILLER_0_249_892 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13199_ VGND VPWR VGND VPWR _07691_ keymem.key_mem\[3\]\[103\] _08698_ _08699_ sky130_fd_sc_hd__a21o_2
XFILLER_0_23_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1049 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19815_ VGND VPWR _00693_ _05317_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_97_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16958_ VPWR VGND VPWR VGND _02603_ _02601_ key[182] _09866_ _03088_ sky130_fd_sc_hd__a22o_2
X_19746_ VGND VPWR _05281_ _05246_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_223_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15909_ VGND VPWR VGND VPWR _11365_ _11273_ _11289_ _11272_ _11288_ sky130_fd_sc_hd__and4_2
X_19677_ VGND VPWR _00628_ _05244_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16889_ VGND VPWR VPWR VGND _02986_ keymem.key_mem\[14\]\[47\] _03025_ _03026_ sky130_fd_sc_hd__mux2_2
XFILLER_0_95_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18628_ VPWR VGND _04496_ enc_block.block_w2_reg\[23\] enc_block.block_w2_reg\[19\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_154_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_133_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_352 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18559_ VPWR VGND _04434_ enc_block.block_w1_reg\[29\] enc_block.block_w2_reg\[21\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_73_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21570_ VGND VPWR _01516_ _06249_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_168_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20521_ VGND VPWR _05692_ _05679_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_6_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_34_219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_28_794 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_248_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23240_ VPWR VGND VPWR VGND _07127_ _04874_ _07125_ enc_block.block_w3_reg\[3\] _07115_
+ _02308_ sky130_fd_sc_hd__a221o_2
X_20452_ VGND VPWR VPWR VGND _05649_ _03550_ keymem.key_mem\[9\]\[109\] _05655_ sky130_fd_sc_hd__mux2_2
XFILLER_0_31_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_403 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23171_ VGND VPWR VPWR VGND _07054_ _07070_ keymem.prev_key1_reg\[119\] _07071_ sky130_fd_sc_hd__mux2_2
X_20383_ VGND VPWR VPWR VGND _05614_ _03295_ keymem.key_mem\[9\]\[76\] _05619_ sky130_fd_sc_hd__mux2_2
XFILLER_0_88_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_1137 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_105_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22122_ VGND VPWR _01773_ _06544_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_109_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_144_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_458 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_112_173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22053_ VGND VPWR _01740_ _06508_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_179_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21004_ VGND VPWR VPWR VGND _05945_ _05054_ keymem.key_mem\[7\]\[110\] _05950_ sky130_fd_sc_hd__mux2_2
XFILLER_0_220_1373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_179_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_103_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25812_ VGND VPWR VPWR VGND clk _02305_ reset_n enc_block.block_w3_reg\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_255_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25743_ keymem.prev_key1_reg\[59\] clk _02236_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22955_ VGND VPWR _02210_ _06940_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_242_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21906_ VPWR VGND keymem.key_mem\[3\]\[20\] _06430_ _06427_ VPWR VGND sky130_fd_sc_hd__and2_2
X_25674_ VGND VPWR VPWR VGND clk _02167_ reset_n keymem.rcon_reg\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_116_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22886_ VGND VPWR VGND VPWR _02184_ _06897_ _06882_ keymem.prev_key1_reg\[7\] sky130_fd_sc_hd__o21a_2
XFILLER_0_151_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_112_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_976 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24625_ VGND VPWR VPWR VGND clk _01118_ reset_n keymem.key_mem\[8\]\[106\] sky130_fd_sc_hd__dfrtp_2
X_21837_ VGND VPWR VPWR VGND _06388_ _03607_ keymem.key_mem\[4\]\[118\] _06391_ sky130_fd_sc_hd__mux2_2
XFILLER_0_52_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_486 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_65_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12570_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[41\] _07724_ keymem.key_mem\[1\]\[41\]
+ _07557_ _08132_ sky130_fd_sc_hd__a22o_2
XFILLER_0_13_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21768_ VGND VPWR _01609_ _06354_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24556_ VGND VPWR VPWR VGND clk _01049_ reset_n keymem.key_mem\[8\]\[37\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_186_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20719_ VGND VPWR VPWR VGND _05794_ _03538_ keymem.key_mem\[8\]\[107\] _05796_ sky130_fd_sc_hd__mux2_2
X_23507_ VGND VPWR VPWR VGND clk _00011_ reset_n result_valid sky130_fd_sc_hd__dfrtp_2
X_24487_ VGND VPWR VPWR VGND clk _00980_ reset_n keymem.key_mem\[9\]\[96\] sky130_fd_sc_hd__dfrtp_2
X_21699_ VGND VPWR _01576_ _06318_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_227_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_266_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14240_ _09639_ _09711_ keymem.prev_key0_reg\[97\] _09709_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_23438_ VGND VPWR _07305_ _04232_ _02328_ _07096_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_262_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14171_ VPWR VGND VGND VPWR _09086_ _09124_ _09140_ _09642_ sky130_fd_sc_hd__nor3_2
XFILLER_0_22_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23369_ VGND VPWR _07244_ enc_block.round_key\[16\] _07243_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_150_257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_260_1142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_123_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13122_ VPWR VGND VPWR VGND _08629_ keymem.key_mem\[5\]\[95\] _08052_ keymem.key_mem\[11\]\[95\]
+ _07902_ _08630_ sky130_fd_sc_hd__a221o_2
X_25108_ VGND VPWR VPWR VGND clk _01601_ reset_n keymem.key_mem\[4\]\[77\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_150_279 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_162_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1295 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_123_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13053_ VGND VPWR enc_block.round_key\[88\] _08567_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17930_ VGND VPWR _00241_ _03884_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25039_ VGND VPWR VPWR VGND clk _01532_ reset_n keymem.key_mem\[4\]\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_218_520 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12004_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[0\] _07536_ _07606_ _07575_ _07607_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_218_542 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17861_ VGND VPWR _00219_ _03837_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_108_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19600_ VGND VPWR VGND VPWR _05202_ keymem.key_mem_we _03444_ _05187_ _00593_ sky130_fd_sc_hd__a31o_2
X_16812_ VGND VPWR VPWR VGND _02884_ keymem.key_mem\[14\]\[40\] _02955_ _02956_ sky130_fd_sc_hd__mux2_2
X_17792_ VGND VPWR VGND VPWR _03732_ keymem.prev_key1_reg\[57\] _03790_ _03789_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_79_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19531_ VGND VPWR VGND VPWR _05166_ keymem.key_mem_we _03150_ _05164_ _00560_ sky130_fd_sc_hd__a31o_2
XFILLER_0_234_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16743_ VPWR VGND VPWR VGND _02892_ _02497_ _02888_ key[162] _02723_ _02893_ sky130_fd_sc_hd__a221o_2
X_13955_ VGND VPWR VGND VPWR _09415_ _09423_ _09381_ _09426_ _09248_ _09427_ sky130_fd_sc_hd__o32a_2
XFILLER_0_233_578 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19462_ VGND VPWR VGND VPWR _05129_ keymem.key_mem_we _02787_ _05121_ _00528_ sky130_fd_sc_hd__a31o_2
X_12906_ VPWR VGND VPWR VGND keymem.key_mem\[8\]\[74\] _07878_ keymem.key_mem\[2\]\[74\]
+ _08131_ _08435_ sky130_fd_sc_hd__a22o_2
XFILLER_0_220_239 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16674_ VGND VPWR VGND VPWR _02815_ _02814_ keymem.prev_key1_reg\[126\] _02828_ sky130_fd_sc_hd__a21o_2
X_13886_ VGND VPWR _09358_ _09357_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18413_ VGND VPWR VPWR VGND enc_block.sword_ctr_inc _07374_ _08945_ _04303_ sky130_fd_sc_hd__or3_2
X_15625_ VGND VPWR VGND VPWR _10633_ _10485_ _10475_ _10459_ _10553_ _11083_ sky130_fd_sc_hd__o32a_2
XFILLER_0_158_335 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12837_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[67\] _07620_ keymem.key_mem\[4\]\[67\]
+ _07636_ _08373_ sky130_fd_sc_hd__a22o_2
X_19393_ VGND VPWR VPWR VGND _04876_ _05089_ keymem.key_mem\[13\]\[127\] _05090_ sky130_fd_sc_hd__mux2_2
XFILLER_0_68_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_29_525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18344_ VPWR VGND VPWR VGND _04241_ _04189_ _04239_ enc_block.block_w0_reg\[24\]
+ _03993_ _00298_ sky130_fd_sc_hd__a221o_2
X_15556_ VPWR VGND VGND VPWR _11015_ _11013_ _11014_ sky130_fd_sc_hd__nand2_2
XFILLER_0_267_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12768_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[60\] _07674_ keymem.key_mem\[12\]\[60\]
+ _07673_ _08311_ sky130_fd_sc_hd__a22o_2
XFILLER_0_29_569 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_210_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1085 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14507_ VGND VPWR VGND VPWR _09080_ _09069_ _09156_ _09083_ _09976_ sky130_fd_sc_hd__o22a_2
XFILLER_0_189_1187 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18275_ VPWR VGND VPWR VGND _04179_ _03970_ _11619_ sky130_fd_sc_hd__or2_2
X_11719_ VGND VPWR result[26] _07423_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15487_ VGND VPWR VGND VPWR _10947_ _10946_ _10943_ _10941_ _10939_ sky130_fd_sc_hd__and4_2
XFILLER_0_71_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12699_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[53\] _08145_ _08248_ _08244_ _08249_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_116_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17226_ VGND VPWR _03330_ _03329_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14438_ VGND VPWR VGND VPWR _09332_ _09323_ _09559_ _09408_ _09907_ sky130_fd_sc_hd__o22a_2
XFILLER_0_4_625 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_64_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17157_ VGND VPWR _03268_ _03267_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_4_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14369_ VGND VPWR VGND VPWR _09140_ _09204_ _09839_ _09167_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_24_285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16108_ VGND VPWR VGND VPWR _11460_ _11218_ _11562_ _11330_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_64_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17088_ VPWR VGND VPWR VGND _09516_ _09854_ _09853_ keymem.prev_key0_reg\[66\] _03206_
+ sky130_fd_sc_hd__or4_2
XFILLER_0_229_818 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16039_ VPWR VGND VGND VPWR _11367_ _11273_ _11227_ _11288_ _11494_ sky130_fd_sc_hd__and4b_2
XFILLER_0_58_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_659 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1100 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_97_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19729_ VGND VPWR _00652_ _05272_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_237_1177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_74_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_205_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22740_ VGND VPWR _02100_ _06835_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_48_801 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22671_ VGND VPWR VPWR VGND _06798_ keymem.key_mem\[0\]\[24\] _02689_ _06807_ sky130_fd_sc_hd__mux2_2
XFILLER_0_181_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21622_ VGND VPWR _01539_ _06278_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24410_ VGND VPWR VPWR VGND clk _00903_ reset_n keymem.key_mem\[9\]\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_34_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25390_ VGND VPWR VPWR VGND clk _01883_ reset_n keymem.key_mem\[2\]\[103\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_191_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_191_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24341_ VGND VPWR VPWR VGND clk _00834_ reset_n keymem.key_mem\[10\]\[78\] sky130_fd_sc_hd__dfrtp_2
X_21553_ VGND VPWR _01508_ _06240_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_69_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_1_Left_403 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20504_ VGND VPWR _01016_ _05683_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24272_ VGND VPWR VPWR VGND clk _00765_ reset_n keymem.key_mem\[10\]\[9\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_140_2_Right_212 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_485 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21484_ VGND VPWR _01475_ _06204_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_69_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_496 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23223_ VPWR VGND VPWR VGND _07111_ block[2] _03958_ enc_block.block_w2_reg\[2\]
+ _03953_ _07112_ sky130_fd_sc_hd__a221o_2
XFILLER_0_209_1257 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_786 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20435_ VGND VPWR VPWR VGND _05638_ _03499_ keymem.key_mem\[9\]\[101\] _05646_ sky130_fd_sc_hd__mux2_2
XFILLER_0_31_723 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_15_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23154_ VGND VPWR VGND VPWR _02288_ _07061_ _07010_ keymem.prev_key1_reg\[111\] sky130_fd_sc_hd__o21a_2
X_20366_ VPWR VGND VGND VPWR _05610_ keymem.key_mem\[9\]\[68\] _05532_ sky130_fd_sc_hd__nand2_2
XFILLER_0_105_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22105_ VGND VPWR _01765_ _06535_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_12_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23085_ VGND VPWR VGND VPWR _07018_ _03379_ _03378_ _03382_ _07011_ sky130_fd_sc_hd__a211o_2
XFILLER_0_105_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20297_ VGND VPWR VPWR VGND _05569_ _02904_ keymem.key_mem\[9\]\[35\] _05574_ sky130_fd_sc_hd__mux2_2
X_22036_ VPWR VGND keymem.key_mem\[3\]\[80\] _06500_ _06484_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_246_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_179_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1192 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_76_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23987_ VGND VPWR VPWR VGND clk _00480_ reset_n keymem.key_mem\[13\]\[108\] sky130_fd_sc_hd__dfrtp_2
X_13740_ VGND VPWR VGND VPWR _09209_ _09160_ _09212_ _09211_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_225_46 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25726_ keymem.prev_key1_reg\[42\] clk _02219_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_225_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22938_ VGND VPWR _02203_ _06930_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_196_953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_57_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_116_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13671_ VPWR VGND VGND VPWR _09069_ _09136_ _09134_ _09132_ _09143_ _09142_ sky130_fd_sc_hd__o221a_2
X_25657_ VGND VPWR VPWR VGND clk _02150_ reset_n keymem.key_mem\[0\]\[114\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_97_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22869_ VGND VPWR VGND VPWR _06886_ _09794_ _03795_ _06884_ _09860_ sky130_fd_sc_hd__a211o_2
XFILLER_0_167_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15410_ VPWR VGND VGND VPWR _10411_ _10495_ _10871_ _10559_ _10510_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_38_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12622_ VPWR VGND VPWR VGND _08178_ keymem.key_mem\[8\]\[46\] _07540_ keymem.key_mem\[1\]\[46\]
+ _07670_ _08179_ sky130_fd_sc_hd__a221o_2
X_24608_ VGND VPWR VPWR VGND clk _01101_ reset_n keymem.key_mem\[8\]\[89\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16390_ VGND VPWR VPWR VGND _11072_ _11089_ keymem.round_ctr_reg\[0\] _02552_ sky130_fd_sc_hd__or3_2
XFILLER_0_167_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1015 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25588_ VGND VPWR VPWR VGND clk _02081_ reset_n keymem.key_mem\[0\]\[45\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_68_1_Left_335 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15341_ VPWR VGND VGND VPWR _10618_ _10803_ _10563_ sky130_fd_sc_hd__nor2_2
X_12553_ VGND VPWR _08116_ _07646_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24539_ VGND VPWR VPWR VGND clk _01032_ reset_n keymem.key_mem\[8\]\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_87_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18060_ VGND VPWR _03981_ _03955_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_120_1_Left_387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15272_ VGND VPWR _10735_ _09932_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_266_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12484_ VPWR VGND VPWR VGND _08053_ keymem.key_mem\[5\]\[33\] _08052_ keymem.key_mem\[3\]\[33\]
+ _07690_ _08054_ sky130_fd_sc_hd__a221o_2
XFILLER_0_87_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17011_ _02757_ _03136_ _03134_ _02758_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_163_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14223_ VGND VPWR VGND VPWR _09033_ _09091_ _09694_ _09056_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_1089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_123_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_149_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1_606 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14154_ VPWR VGND VGND VPWR _09335_ _09327_ _09625_ _09352_ _09293_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_123_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13105_ VGND VPWR enc_block.round_key\[93\] _08614_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_46_1198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_238_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14085_ VGND VPWR VPWR VGND _09248_ _09361_ _09556_ _09464_ _09550_ sky130_fd_sc_hd__o211a_2
X_18962_ VPWR VGND VGND VPWR _04778_ _04797_ _04211_ sky130_fd_sc_hd__nor2_2
XFILLER_0_24_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13036_ VPWR VGND VPWR VGND _08551_ keymem.key_mem\[11\]\[87\] _07781_ keymem.key_mem\[2\]\[87\]
+ _07698_ _08552_ sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_232_Left_499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17913_ VPWR VGND VPWR VGND _03872_ _03871_ keymem.prev_key0_reg\[95\] _03788_ _00236_
+ sky130_fd_sc_hd__a22o_2
X_18893_ VGND VPWR VPWR VGND _04600_ enc_block.block_w2_reg\[14\] _04135_ _04735_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_98_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_158_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_150_2_Left_621 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17844_ VGND VPWR VPWR VGND _03814_ _03825_ keymem.prev_key0_reg\[73\] _03826_ sky130_fd_sc_hd__mux2_2
XFILLER_0_98_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_59_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17775_ VGND VPWR VPWR VGND _03777_ _03062_ keymem.prev_key0_reg\[51\] _03779_ sky130_fd_sc_hd__mux2_2
XFILLER_0_195_1191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14987_ VGND VPWR _10451_ _10412_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_88_200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_238_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19514_ VPWR VGND keymem.key_mem\[12\]\[53\] _05157_ _05128_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16726_ VGND VPWR _02877_ _11543_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13938_ VGND VPWR _09410_ _09409_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_232_1030 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19445_ VPWR VGND keymem.key_mem\[12\]\[21\] _05120_ _05116_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_134_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16657_ VGND VPWR _02812_ _02811_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13869_ VGND VPWR _09341_ _09340_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15608_ VGND VPWR VGND VPWR _10459_ _10569_ _10563_ _10566_ _11066_ sky130_fd_sc_hd__o22a_2
XFILLER_0_31_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19376_ VGND VPWR _00493_ _05078_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_169_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16588_ VPWR VGND VPWR VGND _02745_ keymem.rcon_reg\[3\] sky130_fd_sc_hd__inv_2
XFILLER_0_173_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18327_ VGND VPWR _04226_ enc_block.block_w0_reg\[31\] _04225_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15539_ VPWR VGND VGND VPWR _10534_ _10998_ _10411_ sky130_fd_sc_hd__nor2_2
XFILLER_0_169_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_399 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_60_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18258_ VPWR VGND _04163_ _04079_ enc_block.block_w0_reg\[25\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_245_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_945 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_154_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17209_ VGND VPWR VPWR VGND _03296_ keymem.key_mem\[14\]\[78\] _03314_ _03315_ sky130_fd_sc_hd__mux2_2
XFILLER_0_245_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18189_ VGND VPWR _04100_ _04011_ _04099_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_206_1419 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20220_ VGND VPWR _05532_ _05531_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_163_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_935 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20151_ VGND VPWR _00851_ _05495_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_12_299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_106_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_42_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_2_Left_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20082_ VGND VPWR _00818_ _05459_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_176_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23910_ VGND VPWR VPWR VGND clk _00403_ reset_n keymem.key_mem\[13\]\[31\] sky130_fd_sc_hd__dfrtp_2
X_24890_ VGND VPWR VPWR VGND clk _01383_ reset_n keymem.key_mem\[6\]\[115\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_256_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23841_ VGND VPWR VPWR VGND clk _00334_ reset_n enc_block.block_w1_reg\[26\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_252_1406 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_515 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_174_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_212_526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23772_ VPWR VGND VPWR VGND enc_block.enc_ctrl_reg\[0\] reset_n _00007_ clk sky130_fd_sc_hd__dfstp_2
X_20984_ VGND VPWR _01240_ _05939_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_192_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25511_ VGND VPWR VPWR VGND clk _02004_ reset_n keymem.key_mem\[1\]\[96\] sky130_fd_sc_hd__dfrtp_2
X_22723_ VGND VPWR _02092_ _06826_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_71_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_113_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25442_ VGND VPWR VPWR VGND clk _01935_ reset_n keymem.key_mem\[1\]\[27\] sky130_fd_sc_hd__dfrtp_2
X_22654_ VGND VPWR _06798_ _06784_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_164_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21605_ VGND VPWR _01531_ _06269_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_36_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25373_ VGND VPWR VPWR VGND clk _01866_ reset_n keymem.key_mem\[2\]\[86\] sky130_fd_sc_hd__dfrtp_2
X_22585_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[99\] _06767_ _06766_ _05031_ _02007_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_62_111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24324_ VGND VPWR VPWR VGND clk _00817_ reset_n keymem.key_mem\[10\]\[61\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_263_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21536_ VGND VPWR VPWR VGND _06231_ _03518_ keymem.key_mem\[5\]\[104\] _06232_ sky130_fd_sc_hd__mux2_2
XFILLER_0_145_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_141_2_Right_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21467_ VGND VPWR _01467_ _06195_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24255_ VGND VPWR VPWR VGND clk _00748_ reset_n keymem.key_mem\[11\]\[120\] sky130_fd_sc_hd__dfrtp_2
X_23206_ VGND VPWR _07096_ _07095_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20418_ VGND VPWR VPWR VGND _05627_ _03444_ keymem.key_mem\[9\]\[93\] _05637_ sky130_fd_sc_hd__mux2_2
X_24186_ VGND VPWR VPWR VGND clk _00679_ reset_n keymem.key_mem\[11\]\[51\] sky130_fd_sc_hd__dfrtp_2
X_21398_ VGND VPWR _01434_ _06159_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_120_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_82_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20349_ VGND VPWR VPWR VGND _05591_ _03150_ keymem.key_mem\[9\]\[60\] _05601_ sky130_fd_sc_hd__mux2_2
X_23137_ VGND VPWR VGND VPWR _03529_ _10085_ _03532_ _07050_ sky130_fd_sc_hd__a21o_2
X_23068_ VPWR VGND VPWR VGND _07008_ keymem.prev_key1_reg\[79\] _06926_ sky130_fd_sc_hd__or2_2
XFILLER_0_219_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_200_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14910_ _09165_ _10374_ keymem.prev_key1_reg\[104\] _09238_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_22019_ VGND VPWR _01724_ _06490_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15890_ VGND VPWR VGND VPWR _11278_ _11316_ _11346_ _11345_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_262_459 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_215_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14841_ VPWR VGND VPWR VGND _10299_ _10305_ _10303_ _09470_ _10306_ sky130_fd_sc_hd__or4_2
XFILLER_0_203_526 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17560_ VGND VPWR VGND VPWR _03623_ _02928_ _02877_ key[121] sky130_fd_sc_hd__o21a_2
X_14772_ VGND VPWR VGND VPWR _09582_ _09437_ _09476_ _09366_ _10238_ sky130_fd_sc_hd__o22a_2
X_11984_ VGND VPWR _07587_ _07586_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_153_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16511_ VGND VPWR VPWR VGND _02671_ _02670_ keymem.prev_key0_reg\[120\] keymem.round_ctr_reg\[0\]
+ _02668_ _02669_ sky130_fd_sc_hd__o311ai_2
X_13723_ VGND VPWR VGND VPWR _09194_ _09138_ _09195_ _09136_ sky130_fd_sc_hd__a21oi_2
X_25709_ keymem.prev_key1_reg\[25\] clk _02202_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_17491_ VPWR VGND VGND VPWR _11153_ _03563_ _11152_ sky130_fd_sc_hd__nor2_2
XFILLER_0_85_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19230_ VGND VPWR VPWR VGND _04951_ _04983_ keymem.key_mem\[13\]\[70\] _04984_ sky130_fd_sc_hd__mux2_2
X_16442_ VGND VPWR VPWR VGND _10091_ key[150] keymem.prev_key1_reg\[22\] _02604_ sky130_fd_sc_hd__mux2_2
X_13654_ VPWR VGND VPWR VGND _09031_ _09065_ _09017_ _08957_ _09126_ sky130_fd_sc_hd__or4_2
XFILLER_0_116_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_152 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_195_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19161_ VGND VPWR VPWR VGND _04928_ _04941_ keymem.key_mem\[13\]\[43\] _04942_ sky130_fd_sc_hd__mux2_2
X_12605_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[44\] _08145_ _08163_ _08157_ _08164_
+ sky130_fd_sc_hd__o22a_2
X_16373_ VGND VPWR VGND VPWR _02515_ _02535_ _02536_ _02500_ _02526_ sky130_fd_sc_hd__nor4_2
XFILLER_0_26_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13585_ VGND VPWR _09057_ _09009_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18112_ VPWR VGND VGND VPWR _10917_ _04030_ _08940_ sky130_fd_sc_hd__nor2_2
X_15324_ VPWR VGND VGND VPWR _10536_ _10786_ _10510_ sky130_fd_sc_hd__nor2_2
X_12536_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[38\] _07787_ keymem.key_mem\[2\]\[38\]
+ _07646_ _08101_ sky130_fd_sc_hd__a22o_2
X_19092_ VGND VPWR VGND VPWR _04900_ keymem.key_mem_we _11149_ _04896_ _00387_ sky130_fd_sc_hd__a31o_2
XFILLER_0_42_818 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_48_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18043_ VGND VPWR VGND VPWR _03965_ _07381_ enc_block.sword_ctr_inc enc_block.enc_ctrl_reg\[3\]
+ _07374_ sky130_fd_sc_hd__o211ai_2
X_15255_ VGND VPWR VGND VPWR _10481_ _10587_ _10568_ _10604_ _10718_ sky130_fd_sc_hd__o22a_2
X_12467_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[32\] _07618_ keymem.key_mem\[10\]\[32\]
+ _07742_ _08038_ sky130_fd_sc_hd__a22o_2
XFILLER_0_2_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14206_ VPWR VGND VPWR VGND _09675_ _09676_ _09677_ _09670_ _09674_ sky130_fd_sc_hd__or4b_2
XFILLER_0_111_216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15186_ VPWR VGND VGND VPWR _10480_ _10585_ _10650_ _10649_ _10639_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_160_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12398_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[26\] _07618_ keymem.key_mem\[11\]\[26\]
+ _07761_ _07975_ sky130_fd_sc_hd__a22o_2
XFILLER_0_164_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_111_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_240_Left_507 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14137_ VPWR VGND VGND VPWR _09348_ _09352_ _09608_ _09318_ _09443_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_1_469 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_61_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19994_ VGND VPWR _05413_ _05388_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_226_607 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18945_ VGND VPWR _04781_ enc_block.block_w2_reg\[28\] _04780_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_14068_ VGND VPWR _09540_ _09539_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_59_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13019_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[85\] _07724_ keymem.key_mem\[3\]\[85\]
+ _07843_ _08537_ sky130_fd_sc_hd__a22o_2
XFILLER_0_183_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18876_ VPWR VGND VGND VPWR _04719_ enc_block.block_w1_reg\[4\] enc_block.block_w1_reg\[5\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_207_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17827_ VGND VPWR _03814_ _03673_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_238_1261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_238_1272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_206_397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_171_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17758_ VGND VPWR _00184_ _03769_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_162_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_171_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16709_ VGND VPWR _02862_ _02861_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17689_ VGND VPWR _00162_ _03722_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19428_ VPWR VGND keymem.key_mem\[12\]\[13\] _05111_ _05102_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_130_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19359_ VGND VPWR _05067_ _04876_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_84_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22370_ VGND VPWR VPWR VGND _06669_ _03555_ keymem.key_mem\[2\]\[110\] _06676_ sky130_fd_sc_hd__mux2_2
XFILLER_0_161_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21321_ VGND VPWR _01397_ _06119_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_26_881 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21252_ VGND VPWR _01366_ _06081_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24040_ VGND VPWR VPWR VGND clk _00533_ reset_n keymem.key_mem\[12\]\[33\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_229_401 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20203_ VGND VPWR _00876_ _05522_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21183_ VGND VPWR _01333_ _06045_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_256_231 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1_981 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20134_ VGND VPWR _00843_ _05486_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_256_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_99_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20065_ VGND VPWR _00810_ _05450_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24942_ VGND VPWR VPWR VGND clk _01435_ reset_n keymem.key_mem\[5\]\[39\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24873_ VGND VPWR VPWR VGND clk _01366_ reset_n keymem.key_mem\[6\]\[98\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_172 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23824_ VGND VPWR VPWR VGND clk _00317_ reset_n enc_block.block_w1_reg\[9\] sky130_fd_sc_hd__dfrtp_2
X_23755_ keymem.prev_key0_reg\[111\] clk _00252_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20967_ VGND VPWR VGND VPWR _05930_ keymem.key_mem_we _03435_ _05916_ _01232_ sky130_fd_sc_hd__a31o_2
X_22706_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[45\] _06820_ _06819_ _04945_ _02081_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_177_260 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_137_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_67_269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23686_ keymem.prev_key0_reg\[42\] clk _00183_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_137_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_48_450 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_82_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20898_ VGND VPWR VGND VPWR _05894_ keymem.key_mem_we _03140_ _05893_ _01199_ sky130_fd_sc_hd__a31o_2
XFILLER_0_64_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25425_ VGND VPWR VPWR VGND clk _01918_ reset_n keymem.key_mem\[1\]\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22637_ VGND VPWR _06790_ _06779_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_36_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_442 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_116 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_24_807 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25356_ VGND VPWR VPWR VGND clk _01849_ reset_n keymem.key_mem\[2\]\[69\] sky130_fd_sc_hd__dfrtp_2
X_13370_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[120\] _08216_ keymem.key_mem\[2\]\[120\]
+ _08131_ _08853_ sky130_fd_sc_hd__a22o_2
XFILLER_0_8_580 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_51_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22568_ VGND VPWR _01995_ _06768_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_49_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24307_ VGND VPWR VPWR VGND clk _00800_ reset_n keymem.key_mem\[10\]\[44\] sky130_fd_sc_hd__dfrtp_2
X_12321_ VPWR VGND VPWR VGND _07904_ keymem.key_mem\[11\]\[19\] _07902_ keymem.key_mem\[1\]\[19\]
+ _07901_ _07905_ sky130_fd_sc_hd__a221o_2
XFILLER_0_50_114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21519_ VGND VPWR VPWR VGND _06220_ _03466_ keymem.key_mem\[5\]\[96\] _06223_ sky130_fd_sc_hd__mux2_2
X_25287_ VGND VPWR VPWR VGND clk _01780_ reset_n keymem.key_mem\[2\]\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22499_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[48\] _06737_ _06736_ _04950_ _01956_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_228_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15040_ VGND VPWR _10504_ _10503_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_142_2_Right_214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24238_ VGND VPWR VPWR VGND clk _00731_ reset_n keymem.key_mem\[11\]\[103\] sky130_fd_sc_hd__dfrtp_2
X_12252_ VGND VPWR _07841_ _07693_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_160_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_1282 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_107_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12183_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[10\] _07657_ keymem.key_mem\[9\]\[10\]
+ _07717_ _07776_ sky130_fd_sc_hd__a22o_2
X_24169_ VGND VPWR VPWR VGND clk _00662_ reset_n keymem.key_mem\[11\]\[34\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_82_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16991_ VGND VPWR VGND VPWR _03118_ _11151_ key[185] _03113_ _03117_ sky130_fd_sc_hd__a211o_2
X_15942_ VPWR VGND VPWR VGND _11192_ _11229_ _11207_ _11225_ _11398_ sky130_fd_sc_hd__or4_2
X_18730_ VGND VPWR VGND VPWR _04586_ _04585_ _04587_ _04077_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_159_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1136 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18661_ VPWR VGND VPWR VGND _04525_ block[87] _04487_ enc_block.block_w2_reg\[23\]
+ _04425_ _04526_ sky130_fd_sc_hd__a221o_2
X_15873_ VGND VPWR _11329_ _11328_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_235_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_116_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14824_ VPWR VGND VPWR VGND _10289_ _09368_ _09399_ _09350_ _09898_ _10288_ sky130_fd_sc_hd__o311a_2
X_17612_ VGND VPWR VPWR VGND _09863_ keymem.key_mem\[14\]\[127\] _03668_ _03669_ sky130_fd_sc_hd__mux2_2
X_18592_ VPWR VGND VGND VPWR _04464_ _04401_ _04462_ sky130_fd_sc_hd__nand2_2
XFILLER_0_231_665 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_153_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17543_ VGND VPWR _00130_ _03608_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14755_ _10219_ _10221_ _10218_ _10220_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_93_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11967_ VPWR VGND VPWR VGND _07569_ keymem.key_mem\[10\]\[0\] _07562_ keymem.key_mem\[1\]\[0\]
+ _07558_ _07570_ sky130_fd_sc_hd__a221o_2
XFILLER_0_58_236 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_50_1106 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13706_ VGND VPWR _09178_ _09036_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17474_ VPWR VGND _09533_ _03549_ _03548_ VPWR VGND sky130_fd_sc_hd__and2_2
X_14686_ VGND VPWR VGND VPWR _09110_ _09090_ _10153_ _09116_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_54_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11898_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[20\] dec_new_block\[116\]
+ _07513_ sky130_fd_sc_hd__mux2_2
XFILLER_0_39_461 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16425_ VGND VPWR VGND VPWR _02586_ keymem.round_ctr_reg\[0\] _02587_ _02572_ sky130_fd_sc_hd__nand3_2
X_19213_ VGND VPWR VGND VPWR _04973_ keymem.key_mem_we _03184_ _04968_ _00435_ sky130_fd_sc_hd__a31o_2
X_13637_ VGND VPWR _09109_ _09016_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_55_932 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_128_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19144_ VGND VPWR VGND VPWR _04930_ keymem.key_mem_we _02924_ _04924_ _00409_ sky130_fd_sc_hd__a31o_2
XFILLER_0_143_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16356_ VPWR VGND VPWR VGND _02517_ _02518_ _02519_ _02516_ _02441_ sky130_fd_sc_hd__or4b_2
X_13568_ VGND VPWR _09040_ _09039_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_48_1002 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_143_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15307_ VGND VPWR VGND VPWR _10769_ _10633_ _10554_ _10540_ sky130_fd_sc_hd__o21a_2
XFILLER_0_246_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12519_ VGND VPWR enc_block.round_key\[36\] _08085_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19075_ VPWR VGND keymem.key_mem\[13\]\[8\] _04891_ _04887_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16287_ VGND VPWR VGND VPWR _02451_ _11432_ _11396_ _11365_ _11348_ _11224_ sky130_fd_sc_hd__a32o_2
XFILLER_0_2_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13499_ VGND VPWR _08971_ _08970_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_207_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18026_ VGND VPWR VGND VPWR _07374_ _07381_ _03947_ _03948_ sky130_fd_sc_hd__a21o_2
X_15238_ VPWR VGND VGND VPWR _10535_ _10701_ _10521_ sky130_fd_sc_hd__nor2_2
XFILLER_0_41_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_164_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_670 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_125_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15169_ VGND VPWR _10633_ _10623_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_61_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_765 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_142_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_254_724 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19977_ VGND VPWR _00768_ _05404_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18928_ VPWR VGND VGND VPWR _04765_ _04766_ _04478_ sky130_fd_sc_hd__nor2_2
XFILLER_0_66_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_242_919 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_253_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18859_ VPWR VGND VGND VPWR _04704_ _04627_ _04702_ sky130_fd_sc_hd__nand2_2
XFILLER_0_235_982 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_145_1_Left_412 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_96_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21870_ VGND VPWR VGND VPWR _06410_ keymem.key_mem_we _09992_ _06404_ _01655_ sky130_fd_sc_hd__a31o_2
XFILLER_0_89_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_974 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_72_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_132_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20821_ VPWR VGND keymem.key_mem\[7\]\[24\] _05853_ _05844_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_49_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_82_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_136_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23540_ VGND VPWR VPWR VGND clk _00041_ reset_n keymem.key_mem\[14\]\[29\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20752_ VGND VPWR VPWR VGND _05805_ _03640_ keymem.key_mem\[8\]\[123\] _05813_ sky130_fd_sc_hd__mux2_2
X_23471_ VGND VPWR _07334_ _04258_ _02332_ _07115_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_20683_ VGND VPWR VPWR VGND _05772_ _03417_ keymem.key_mem\[8\]\[90\] _05777_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_431 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25210_ VGND VPWR VPWR VGND clk _01703_ reset_n keymem.key_mem\[3\]\[51\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_18_667 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_1_Right_670 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_134_116 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22422_ VGND VPWR _01913_ _06704_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_134_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1174 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_60_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25141_ VGND VPWR VPWR VGND clk _01634_ reset_n keymem.key_mem\[4\]\[110\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22353_ VGND VPWR VPWR VGND _06658_ _03506_ keymem.key_mem\[2\]\[102\] _06667_ sky130_fd_sc_hd__mux2_2
XFILLER_0_5_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21304_ VGND VPWR _01391_ _06108_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_60_467 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22284_ VGND VPWR VPWR VGND _06622_ _03234_ keymem.key_mem\[2\]\[69\] _06631_ sky130_fd_sc_hd__mux2_2
X_25072_ VGND VPWR VPWR VGND clk _01565_ reset_n keymem.key_mem\[4\]\[41\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1046 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_361 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_83_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_143_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21235_ VGND VPWR _01358_ _06072_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24023_ VGND VPWR VPWR VGND clk _00516_ reset_n keymem.key_mem\[12\]\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_130_388 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_44_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_223_1382 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_2_Left_579 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21166_ VGND VPWR _01325_ _06036_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20117_ VGND VPWR _00835_ _05477_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21097_ VGND VPWR _01292_ _06000_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_77_1_Left_344 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_254_1309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_176_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_1231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20048_ VGND VPWR _00802_ _05441_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24925_ VGND VPWR VPWR VGND clk _01418_ reset_n keymem.key_mem\[5\]\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_260_749 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12870_ VGND VPWR VGND VPWR _08403_ _07580_ keymem.key_mem\[12\]\[70\] _08400_ _08402_
+ sky130_fd_sc_hd__a211o_2
X_24856_ VGND VPWR VPWR VGND clk _01349_ reset_n keymem.key_mem\[6\]\[81\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_154_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11821_ VGND VPWR result[77] _07474_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23807_ VGND VPWR VPWR VGND clk _00300_ reset_n enc_block.block_w0_reg\[26\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_90_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24787_ VGND VPWR VPWR VGND clk _01280_ reset_n keymem.key_mem\[6\]\[12\] sky130_fd_sc_hd__dfrtp_2
X_21999_ VPWR VGND keymem.key_mem\[3\]\[63\] _06480_ _06469_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_201_849 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_197_377 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_154_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14540_ VPWR VGND VGND VPWR _09222_ _10008_ _09113_ sky130_fd_sc_hd__nor2_2
X_11752_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[11\] dec_new_block\[43\]
+ _07440_ sky130_fd_sc_hd__mux2_2
XFILLER_0_90_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23738_ keymem.prev_key0_reg\[94\] clk _00235_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_409 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_51_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14471_ VGND VPWR VPWR VGND _09940_ _09020_ _09694_ _09939_ _09181_ sky130_fd_sc_hd__o31a_2
X_11683_ VGND VPWR result[8] _07405_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_165_252 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23669_ keymem.prev_key0_reg\[25\] clk _00166_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_113_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16210_ VGND VPWR VGND VPWR _11482_ _11284_ _02375_ _11306_ sky130_fd_sc_hd__a21oi_2
X_25408_ VGND VPWR VPWR VGND clk _01901_ reset_n keymem.key_mem\[2\]\[121\] sky130_fd_sc_hd__dfrtp_2
X_13422_ VPWR VGND VPWR VGND _08899_ keymem.key_mem\[6\]\[125\] _07711_ keymem.key_mem\[2\]\[125\]
+ _07647_ _08900_ sky130_fd_sc_hd__a221o_2
XFILLER_0_37_976 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17190_ VGND VPWR _00088_ _03297_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16141_ VPWR VGND VGND VPWR _11283_ _11595_ _11284_ sky130_fd_sc_hd__nor2_2
X_25339_ VGND VPWR VPWR VGND clk _01832_ reset_n keymem.key_mem\[2\]\[52\] sky130_fd_sc_hd__dfrtp_2
X_13353_ VGND VPWR VGND VPWR _07842_ keymem.key_mem\[9\]\[118\] _08833_ _08835_ _08838_
+ _08837_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_23_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1282 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12304_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[18\] _07608_ keymem.key_mem\[1\]\[18\]
+ _07556_ _07889_ sky130_fd_sc_hd__a22o_2
XFILLER_0_161_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16072_ VGND VPWR _11527_ _11327_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_23_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_51_478 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13284_ VGND VPWR VGND VPWR _08776_ _07968_ keymem.key_mem\[9\]\[111\] _08773_ _08775_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_165_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_32_670 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15023_ VGND VPWR VGND VPWR _10487_ _10445_ _10430_ _10457_ _10443_ sky130_fd_sc_hd__and4_2
X_19900_ VGND VPWR VPWR VGND _05361_ keymem.key_mem\[11\]\[106\] _03533_ _05362_ sky130_fd_sc_hd__mux2_2
XFILLER_0_161_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_143_2_Right_215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_62_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12235_ VPWR VGND VPWR VGND _07824_ keymem.key_mem\[3\]\[13\] _07602_ keymem.key_mem\[9\]\[13\]
+ _07591_ _07825_ sky130_fd_sc_hd__a221o_2
XFILLER_0_258_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19831_ VGND VPWR _00701_ _05325_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_20_887 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12166_ VGND VPWR _07761_ _07599_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_202_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_236_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19762_ VGND VPWR _00668_ _05289_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_194_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12097_ VGND VPWR _07695_ _07694_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_208_459 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16974_ VPWR VGND VPWR VGND _03102_ key[56] _09719_ sky130_fd_sc_hd__or2_2
XFILLER_0_224_919 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18713_ _04570_ _04572_ _04560_ _04571_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_15925_ VGND VPWR VGND VPWR _11380_ _11253_ _11379_ _11275_ _11377_ _11381_ sky130_fd_sc_hd__o32a_2
X_19693_ VGND VPWR _00635_ _05253_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_194_1278 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15856_ VPWR VGND VPWR VGND _11265_ _11248_ _11243_ _11232_ _11312_ sky130_fd_sc_hd__or4_2
X_18644_ VGND VPWR _04511_ enc_block.round_key\[85\] _04510_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_172_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14807_ VGND VPWR VGND VPWR _10261_ _10243_ _10273_ keymem.prev_key1_reg\[102\] sky130_fd_sc_hd__a21oi_2
XFILLER_0_59_523 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15787_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[17\] _08955_ _11243_ _08942_ _11177_
+ _11178_ sky130_fd_sc_hd__a32oi_2
X_18575_ VPWR VGND VPWR VGND _04448_ block[78] _04351_ enc_block.block_w3_reg\[14\]
+ _03954_ _04449_ sky130_fd_sc_hd__a221o_2
XFILLER_0_133_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12999_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[83\] _07667_ keymem.key_mem\[8\]\[83\]
+ _07903_ _08519_ sky130_fd_sc_hd__a22o_2
XFILLER_0_15_1001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14738_ _10202_ _10204_ _10201_ _10203_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_17526_ VGND VPWR VPWR VGND _03593_ keymem.key_mem\[14\]\[116\] _03592_ _03594_ sky130_fd_sc_hd__mux2_2
XFILLER_0_47_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_15_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_79 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_46_217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17457_ VGND VPWR VPWR VGND _03534_ keymem.key_mem\[14\]\[106\] _03533_ _03535_ sky130_fd_sc_hd__mux2_2
X_14669_ VGND VPWR VGND VPWR _09472_ _09425_ _09478_ _09391_ _09383_ _10136_ sky130_fd_sc_hd__o41a_2
XPHY_EDGE_ROW_91_2_Left_562 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_200_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_15_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16408_ VPWR VGND VGND VPWR _11482_ _11386_ _11379_ _11422_ _02570_ _02569_ sky130_fd_sc_hd__o221a_2
XFILLER_0_89_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17388_ VGND VPWR VPWR VGND _03467_ keymem.key_mem\[14\]\[97\] _03474_ _03475_ sky130_fd_sc_hd__mux2_2
XFILLER_0_109_190 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16339_ VGND VPWR VGND VPWR _11218_ _11302_ _11204_ _11313_ _02502_ sky130_fd_sc_hd__o22a_2
X_19127_ VGND VPWR VGND VPWR _04919_ keymem.key_mem_we _02862_ _04908_ _00403_ sky130_fd_sc_hd__a31o_2
X_19058_ VGND VPWR VGND VPWR _04881_ keymem.key_mem_we _09537_ _04878_ _00372_ sky130_fd_sc_hd__a31o_2
XFILLER_0_112_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_2_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18009_ VGND VPWR VGND VPWR _03938_ _03937_ _03675_ _03659_ sky130_fd_sc_hd__and3b_2
XFILLER_0_168_54 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21020_ VGND VPWR _01257_ _05958_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_168_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_584 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_22_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_263_Right_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22971_ VGND VPWR VPWR VGND _02950_ _02948_ _06950_ _06881_ _02953_ sky130_fd_sc_hd__o211a_2
XFILLER_0_39_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24710_ VGND VPWR VPWR VGND clk _01203_ reset_n keymem.key_mem\[7\]\[63\] sky130_fd_sc_hd__dfrtp_2
X_21922_ VGND VPWR VGND VPWR _06438_ keymem.key_mem_we _02765_ _06432_ _01679_ sky130_fd_sc_hd__a31o_2
X_25690_ keymem.prev_key1_reg\[6\] clk _02183_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_184_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24641_ VGND VPWR VPWR VGND clk _01134_ reset_n keymem.key_mem\[8\]\[122\] sky130_fd_sc_hd__dfrtp_2
X_21853_ VGND VPWR VPWR VGND _06262_ _03661_ keymem.key_mem\[4\]\[126\] _06399_ sky130_fd_sc_hd__mux2_2
XFILLER_0_77_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_136_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20804_ VGND VPWR VGND VPWR _05843_ keymem.key_mem_we _11447_ _05838_ _01156_ sky130_fd_sc_hd__a31o_2
XFILLER_0_38_718 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24572_ VGND VPWR VPWR VGND clk _01065_ reset_n keymem.key_mem\[8\]\[53\] sky130_fd_sc_hd__dfrtp_2
X_21784_ VGND VPWR VPWR VGND _06355_ _03443_ keymem.key_mem\[4\]\[93\] _06363_ sky130_fd_sc_hd__mux2_2
XFILLER_0_72_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23523_ VGND VPWR VPWR VGND clk _00024_ reset_n keymem.key_mem\[14\]\[12\] sky130_fd_sc_hd__dfrtp_2
X_20735_ VGND VPWR VPWR VGND _05794_ _03585_ keymem.key_mem\[8\]\[115\] _05804_ sky130_fd_sc_hd__mux2_2
XFILLER_0_203_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_19_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23454_ VPWR VGND VGND VPWR _07319_ enc_block.block_w3_reg\[25\] enc_block.block_w1_reg\[10\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_68_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20666_ VGND VPWR VPWR VGND _05761_ _03346_ keymem.key_mem\[8\]\[82\] _05768_ sky130_fd_sc_hd__mux2_2
XFILLER_0_188_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22405_ VGND VPWR VPWR VGND _06553_ _03668_ keymem.key_mem\[2\]\[127\] _06694_ sky130_fd_sc_hd__mux2_2
X_23385_ VPWR VGND VGND VPWR _07258_ _07184_ _07257_ sky130_fd_sc_hd__nand2_2
X_20597_ VGND VPWR VPWR VGND _05725_ _03046_ keymem.key_mem\[8\]\[49\] _05732_ sky130_fd_sc_hd__mux2_2
XFILLER_0_6_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25124_ VGND VPWR VPWR VGND clk _01617_ reset_n keymem.key_mem\[4\]\[93\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_225_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22336_ VGND VPWR _06658_ _06552_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_260_1346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_130_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25055_ VGND VPWR VPWR VGND clk _01548_ reset_n keymem.key_mem\[4\]\[24\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_108_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22267_ VGND VPWR _06622_ _06552_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12020_ VGND VPWR _07622_ _07586_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24006_ VGND VPWR VPWR VGND clk _00499_ reset_n keymem.key_mem\[13\]\[127\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_40_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21218_ VGND VPWR _01350_ _06063_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22198_ VGND VPWR VPWR VGND _06578_ _02786_ keymem.key_mem\[2\]\[28\] _06586_ sky130_fd_sc_hd__mux2_2
XFILLER_0_143_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_724 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1231 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21149_ VGND VPWR _01317_ _06027_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_217_234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_206_919 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_79_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13971_ VGND VPWR _09443_ _09442_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15710_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[18\] _08989_ _11166_ _08983_ _11164_
+ _11165_ sky130_fd_sc_hd__a32oi_2
X_12922_ VGND VPWR _08449_ _07534_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24908_ VGND VPWR VPWR VGND clk _01401_ reset_n keymem.key_mem\[5\]\[5\] sky130_fd_sc_hd__dfrtp_2
X_16690_ VGND VPWR keymem.rcon_logic.tmp_rcon\[0\] _02841_ _02843_ _02842_ VPWR VGND
+ sky130_fd_sc_hd__o21ai_2
X_15641_ VGND VPWR _11099_ _11098_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_154_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24839_ VGND VPWR VPWR VGND clk _01332_ reset_n keymem.key_mem\[6\]\[64\] sky130_fd_sc_hd__dfrtp_2
X_12853_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[69\] _07744_ keymem.key_mem\[4\]\[69\]
+ _07636_ _08387_ sky130_fd_sc_hd__a22o_2
XFILLER_0_115_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11804_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[5\] dec_new_block\[69\]
+ _07466_ sky130_fd_sc_hd__mux2_2
X_18360_ VPWR VGND VGND VPWR _04256_ _04004_ _09790_ sky130_fd_sc_hd__nand2_2
XFILLER_0_154_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15572_ _10168_ _11031_ keymem.prev_key1_reg\[109\] _10184_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_12784_ VGND VPWR VGND VPWR _08325_ _07648_ keymem.key_mem\[2\]\[62\] _08324_ _07896_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_90_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17311_ VGND VPWR VGND VPWR key[89] _08937_ _03405_ _03404_ _03406_ sky130_fd_sc_hd__o22a_2
XFILLER_0_16_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14523_ VGND VPWR _09992_ _09991_ VPWR VGND sky130_fd_sc_hd__buf_1
X_11735_ VGND VPWR result[34] _07431_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18291_ VPWR VGND _04193_ enc_block.block_w1_reg\[23\] enc_block.block_w1_reg\[19\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_113_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_548 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_12_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17242_ VGND VPWR VPWR VGND _11624_ _11622_ keymem.prev_key0_reg\[82\] _03344_ sky130_fd_sc_hd__or3_2
X_14454_ VGND VPWR VGND VPWR _09896_ _09922_ _09923_ _09887_ _09909_ sky130_fd_sc_hd__nor4_2
XFILLER_0_260_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11666_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[0\] dec_new_block\[0\]
+ _07397_ sky130_fd_sc_hd__mux2_2
XFILLER_0_86_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13405_ VGND VPWR enc_block.round_key\[123\] _08884_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17173_ VPWR VGND _10894_ _03282_ _10895_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_98_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14385_ VPWR VGND _09855_ keymem.prev_key0_reg\[66\] keymem.prev_key0_reg\[34\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
X_16124_ VPWR VGND VGND VPWR _11397_ _11578_ _11527_ sky130_fd_sc_hd__nor2_2
XFILLER_0_52_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13336_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[117\] _07788_ keymem.key_mem\[4\]\[117\]
+ _07914_ _08822_ sky130_fd_sc_hd__a22o_2
XFILLER_0_45_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_489 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_126_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_161_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16055_ VGND VPWR VGND VPWR _11509_ _11323_ _11409_ _11230_ _11510_ sky130_fd_sc_hd__a31o_2
XFILLER_0_45_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13267_ VGND VPWR enc_block.round_key\[109\] _08760_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_126_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_808 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_161_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15006_ VGND VPWR VGND VPWR _10462_ _10465_ _10469_ _10467_ _10470_ sky130_fd_sc_hd__o22a_2
XPHY_EDGE_ROW_144_2_Right_216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12218_ VGND VPWR _07809_ _07631_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_23_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_259_1017 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13198_ VPWR VGND VPWR VGND keymem.key_mem\[8\]\[103\] _07878_ keymem.key_mem\[2\]\[103\]
+ _07733_ _08698_ sky130_fd_sc_hd__a22o_2
XFILLER_0_62_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19814_ VGND VPWR VPWR VGND _05314_ keymem.key_mem\[11\]\[65\] _03202_ _05317_ sky130_fd_sc_hd__mux2_2
XFILLER_0_138_46 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12149_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[7\] _07744_ keymem.key_mem\[11\]\[7\]
+ _07631_ _07745_ sky130_fd_sc_hd__a22o_2
XFILLER_0_208_234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_97_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19745_ VGND VPWR _00660_ _05280_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16957_ VPWR VGND VPWR VGND _03087_ key[54] _09795_ sky130_fd_sc_hd__or2_2
XFILLER_0_263_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15908_ VPWR VGND VPWR VGND _11342_ _11363_ _11354_ _11322_ _11364_ sky130_fd_sc_hd__or4_2
XFILLER_0_56_1123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19676_ VGND VPWR VPWR VGND _05243_ keymem.key_mem\[11\]\[0\] _09537_ _05244_ sky130_fd_sc_hd__mux2_2
X_16888_ VGND VPWR _03025_ _03024_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_232_760 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18627_ VPWR VGND VPWR VGND _04495_ _04459_ _04494_ enc_block.block_w1_reg\[19\]
+ _04424_ _00327_ sky130_fd_sc_hd__a221o_2
XFILLER_0_188_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_172_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15839_ VGND VPWR _11295_ _11294_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_133_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_172_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18558_ VPWR VGND VPWR VGND _04433_ _04291_ _04432_ enc_block.block_w1_reg\[12\]
+ _04424_ _00320_ sky130_fd_sc_hd__a221o_2
XFILLER_0_133_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_537 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17509_ VPWR VGND VGND VPWR _03578_ _03579_ keylen sky130_fd_sc_hd__nor2_2
X_18489_ VPWR VGND VPWR VGND _04371_ _04291_ _04370_ enc_block.block_w1_reg\[5\] _04317_
+ _00313_ sky130_fd_sc_hd__a221o_2
XFILLER_0_30_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_690 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20520_ VGND VPWR _01024_ _05691_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_34_209 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_184_391 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20451_ VGND VPWR _00992_ _05654_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_248_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_166_1166 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_31_916 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23170_ VGND VPWR VGND VPWR _03609_ _10085_ _03612_ _07070_ sky130_fd_sc_hd__a21o_2
X_20382_ VGND VPWR _05618_ _03287_ _00959_ _05532_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_144_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_990 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_88_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22121_ VGND VPWR VPWR VGND _06538_ _05077_ keymem.key_mem\[3\]\[121\] _06544_ sky130_fd_sc_hd__mux2_2
XFILLER_0_2_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_105_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_247_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22052_ VGND VPWR VPWR VGND _06494_ _05013_ keymem.key_mem\[3\]\[88\] _06508_ sky130_fd_sc_hd__mux2_2
XFILLER_0_80_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_178 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_140_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_255_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21003_ VGND VPWR _01249_ _05949_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_41_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25811_ keymem.prev_key1_reg\[127\] clk _02304_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_255_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25742_ keymem.prev_key1_reg\[58\] clk _02235_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22954_ VGND VPWR VPWR VGND _06914_ _06939_ keymem.prev_key1_reg\[33\] _06940_ sky130_fd_sc_hd__mux2_2
X_21905_ VGND VPWR VGND VPWR _06429_ keymem.key_mem_we _02410_ _06420_ _01671_ sky130_fd_sc_hd__a31o_2
XFILLER_0_218_1281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_190_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25673_ VGND VPWR VPWR VGND clk _02166_ reset_n keymem.rcon_reg\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_155_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22885_ VGND VPWR VGND VPWR _06897_ _10324_ _10321_ _06884_ _10368_ sky130_fd_sc_hd__a211o_2
XFILLER_0_214_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24624_ VGND VPWR VPWR VGND clk _01117_ reset_n keymem.key_mem\[8\]\[105\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_151_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21836_ VGND VPWR _01641_ _06390_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_65_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_112_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24555_ VGND VPWR VPWR VGND clk _01048_ reset_n keymem.key_mem\[8\]\[36\] sky130_fd_sc_hd__dfrtp_2
X_21767_ VGND VPWR VPWR VGND _06344_ _03374_ keymem.key_mem\[4\]\[85\] _06354_ sky130_fd_sc_hd__mux2_2
XFILLER_0_231_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23506_ VGND VPWR _02336_ _07365_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20718_ VGND VPWR _01118_ _05795_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_19_773 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24486_ VGND VPWR VPWR VGND clk _00979_ reset_n keymem.key_mem\[9\]\[95\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_266_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21698_ VGND VPWR VPWR VGND _06308_ _03075_ keymem.key_mem\[4\]\[52\] _06318_ sky130_fd_sc_hd__mux2_2
XFILLER_0_46_570 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23437_ VGND VPWR VGND VPWR _07304_ _04149_ _07095_ _07305_ enc_block.block_w3_reg\[23\]
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_92_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_266_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20649_ VPWR VGND VGND VPWR _05676_ _05759_ keymem.key_mem\[8\]\[74\] sky130_fd_sc_hd__nor2_2
XFILLER_0_135_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14170_ VPWR VGND VGND VPWR _09011_ _09185_ _09157_ _09641_ sky130_fd_sc_hd__nor3_2
X_23368_ VPWR VGND VPWR VGND _07242_ block[16] _04139_ enc_block.block_w0_reg\[16\]
+ _03953_ _07243_ sky130_fd_sc_hd__a221o_2
XFILLER_0_22_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13121_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[95\] _07694_ keymem.key_mem\[12\]\[95\]
+ _07673_ _08629_ sky130_fd_sc_hd__a22o_2
X_25107_ VGND VPWR VPWR VGND clk _01600_ reset_n keymem.key_mem\[4\]\[76\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22319_ VGND VPWR _01865_ _06649_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23299_ VPWR VGND VPWR VGND _07180_ block[9] _04139_ enc_block.block_w1_reg\[9\]
+ _03953_ _07181_ sky130_fd_sc_hd__a221o_2
XFILLER_0_123_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_30_971 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13052_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[88\] _08449_ _08566_ _08562_ _08567_
+ sky130_fd_sc_hd__o22a_2
X_25038_ VGND VPWR VPWR VGND clk _01531_ reset_n keymem.key_mem\[4\]\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_123_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12003_ VGND VPWR VGND VPWR _07606_ _07580_ keymem.key_mem\[12\]\[0\] _07589_ _07605_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_44_1093 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17860_ VGND VPWR VPWR VGND _03836_ _03835_ keymem.prev_key0_reg\[78\] _03837_ sky130_fd_sc_hd__mux2_2
XFILLER_0_79_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16811_ VGND VPWR VGND VPWR _02955_ _02953_ _02950_ _02948_ _02954_ sky130_fd_sc_hd__o211ai_2
X_17791_ VGND VPWR _03789_ _03281_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_260_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_79_1189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19530_ VPWR VGND keymem.key_mem\[12\]\[60\] _05166_ _05158_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13954_ VGND VPWR _09426_ _09425_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16742_ VGND VPWR VPWR VGND _02889_ _09855_ _02892_ _02891_ _02890_ sky130_fd_sc_hd__o211a_2
XFILLER_0_17_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12905_ VGND VPWR VGND VPWR _07800_ keymem.key_mem\[1\]\[74\] _08431_ _08433_ _08434_
+ _08243_ sky130_fd_sc_hd__a2111o_2
X_19461_ VPWR VGND keymem.key_mem\[12\]\[28\] _05129_ _05128_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_220_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16673_ VGND VPWR VPWR VGND _11109_ _02826_ key[30] _02827_ sky130_fd_sc_hd__mux2_2
X_13885_ VGND VPWR _09357_ _09356_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_124_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_213_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18412_ VPWR VGND VPWR VGND _04302_ _04291_ _04300_ enc_block.block_w0_reg\[31\]
+ _03993_ _00305_ sky130_fd_sc_hd__a221o_2
X_15624_ VGND VPWR VGND VPWR _10646_ _10520_ _10618_ _10751_ _11082_ sky130_fd_sc_hd__o22a_2
X_12836_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[67\] _07587_ keymem.key_mem\[3\]\[67\]
+ _07603_ _08372_ sky130_fd_sc_hd__a22o_2
XFILLER_0_75_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19392_ VPWR VGND keymem.key_mem_we _05089_ _03668_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_57_835 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_130_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15555_ VGND VPWR VGND VPWR _10459_ _10480_ _10583_ _11014_ sky130_fd_sc_hd__a21o_2
XFILLER_0_29_537 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18343_ VPWR VGND VGND VPWR _04240_ _04241_ _04190_ sky130_fd_sc_hd__nor2_2
XFILLER_0_210_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12767_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[60\] _07838_ keymem.key_mem\[2\]\[60\]
+ _07816_ _08310_ sky130_fd_sc_hd__a22o_2
XFILLER_0_83_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14506_ VPWR VGND VGND VPWR _09116_ _09109_ _09110_ _09058_ _09975_ _09974_ sky130_fd_sc_hd__o221a_2
XFILLER_0_12_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18274_ VPWR VGND _04178_ _04177_ enc_block.round_key\[114\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_11718_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[26\] dec_new_block\[26\]
+ _07423_ sky130_fd_sc_hd__mux2_2
XFILLER_0_210_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15486_ VGND VPWR VGND VPWR _10946_ _10945_ _10791_ _10790_ _10783_ sky130_fd_sc_hd__and4_2
XFILLER_0_51_1097 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12698_ VGND VPWR VGND VPWR _08248_ _08008_ keymem.key_mem\[2\]\[53\] _08245_ _08247_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_71_326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14437_ VGND VPWR VGND VPWR _09480_ _09476_ _09487_ _09444_ _09906_ sky130_fd_sc_hd__o22a_2
XFILLER_0_71_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17225_ VGND VPWR VGND VPWR _11151_ key[208] _03328_ _03329_ sky130_fd_sc_hd__a21o_2
X_11649_ VGND VPWR _07386_ _07385_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_181_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_126_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_109_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17156_ VGND VPWR VGND VPWR _08930_ key[201] _03266_ _03267_ sky130_fd_sc_hd__a21o_2
X_14368_ VPWR VGND VPWR VGND _09834_ _09213_ _09836_ _09837_ _09838_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_68_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_64_1425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_154_1_Left_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_52_584 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_735 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16107_ VGND VPWR _11561_ keymem.prev_key0_reg\[18\] _11560_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13319_ VGND VPWR VGND VPWR _07780_ keymem.key_mem\[5\]\[115\] _08804_ _08806_ _08807_
+ _08736_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_40_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17087_ VGND VPWR VPWR VGND _09854_ _09853_ _03205_ _08936_ keymem.prev_key0_reg\[66\]
+ sky130_fd_sc_hd__o211a_2
X_14299_ VGND VPWR VPWR VGND _09764_ _09768_ _09454_ _09769_ sky130_fd_sc_hd__or3_2
XFILLER_0_64_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16038_ VPWR VGND VGND VPWR _11482_ _11493_ _11372_ sky130_fd_sc_hd__nor2_2
XFILLER_0_149_67 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_58_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_145_2_Right_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1060 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_671 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_165_11 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17989_ VGND VPWR _00260_ _03924_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_58_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_321 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_263_181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_74_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19728_ VGND VPWR VPWR VGND _05270_ keymem.key_mem\[11\]\[24\] _02689_ _05272_ sky130_fd_sc_hd__mux2_2
XFILLER_0_165_66 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_251_354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_233_1009 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_205_760 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19659_ VGND VPWR _00621_ _05233_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_204_292 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_48_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22670_ VGND VPWR _02059_ _06806_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_90_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1192 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21621_ VGND VPWR VPWR VGND _06275_ _11148_ keymem.key_mem\[4\]\[15\] _06278_ sky130_fd_sc_hd__mux2_2
XFILLER_0_176_166 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_34_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_879 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_69_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_117_2_Left_588 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24340_ VGND VPWR VPWR VGND clk _00833_ reset_n keymem.key_mem\[10\]\[77\] sky130_fd_sc_hd__dfrtp_2
X_21552_ VGND VPWR VPWR VGND _06231_ _03567_ keymem.key_mem\[5\]\[112\] _06240_ sky130_fd_sc_hd__mux2_2
XFILLER_0_1_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_69_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20503_ VGND VPWR VPWR VGND _05680_ _10098_ keymem.key_mem\[8\]\[4\] _05683_ sky130_fd_sc_hd__mux2_2
X_24271_ VGND VPWR VPWR VGND clk _00764_ reset_n keymem.key_mem\[10\]\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_1_Left_353 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21483_ VGND VPWR VPWR VGND _06196_ _03321_ keymem.key_mem\[5\]\[79\] _06204_ sky130_fd_sc_hd__mux2_2
X_23222_ VPWR VGND VGND VPWR _07110_ _07111_ _04382_ sky130_fd_sc_hd__nor2_2
X_20434_ VGND VPWR _00984_ _05645_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_15_264 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_798 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_222_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23153_ VGND VPWR VGND VPWR _07061_ _03557_ _03020_ _06924_ _03559_ sky130_fd_sc_hd__a211o_2
X_20365_ VGND VPWR _00951_ _05609_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_105_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22104_ VGND VPWR VPWR VGND _06527_ _05060_ keymem.key_mem\[3\]\[113\] _06535_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_179_2_Left_650 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_971 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_144_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_278 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23084_ VGND VPWR VGND VPWR _02262_ _07017_ _07010_ keymem.prev_key1_reg\[85\] sky130_fd_sc_hd__o21a_2
XFILLER_0_100_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20296_ VGND VPWR _00918_ _05573_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_219_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22035_ VGND VPWR VGND VPWR _06499_ keymem.key_mem_we _03322_ _06498_ _01731_ sky130_fd_sc_hd__a31o_2
XFILLER_0_179_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23986_ VGND VPWR VPWR VGND clk _00479_ reset_n keymem.key_mem\[13\]\[107\] sky130_fd_sc_hd__dfrtp_2
X_25725_ keymem.prev_key1_reg\[41\] clk _02218_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22937_ VGND VPWR VPWR VGND _06914_ _06929_ keymem.prev_key1_reg\[26\] _06930_ sky130_fd_sc_hd__mux2_2
XFILLER_0_196_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_225_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13670_ VGND VPWR VGND VPWR _09138_ _09125_ _09141_ _09140_ _09142_ sky130_fd_sc_hd__o22a_2
X_25656_ VGND VPWR VPWR VGND clk _02149_ reset_n keymem.key_mem\[0\]\[113\] sky130_fd_sc_hd__dfrtp_2
X_22868_ VGND VPWR VGND VPWR _02178_ _06885_ _06882_ keymem.prev_key1_reg\[1\] sky130_fd_sc_hd__o21a_2
XFILLER_0_38_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_116_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24607_ VGND VPWR VPWR VGND clk _01100_ reset_n keymem.key_mem\[8\]\[88\] sky130_fd_sc_hd__dfrtp_2
X_12621_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[46\] _07602_ keymem.key_mem\[10\]\[46\]
+ _07560_ _08178_ sky130_fd_sc_hd__a22o_2
XFILLER_0_196_987 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_796 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21819_ VGND VPWR _01633_ _06381_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_13_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25587_ VGND VPWR VPWR VGND clk _02080_ reset_n keymem.key_mem\[0\]\[44\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_249_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22799_ VGND VPWR _06857_ _03733_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15340_ VPWR VGND VGND VPWR _10480_ _10528_ _10802_ _10633_ _10612_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_249_1027 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_87_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12552_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[40\] _07691_ keymem.key_mem\[11\]\[40\]
+ _07912_ _08115_ sky130_fd_sc_hd__a22o_2
X_24538_ VGND VPWR VPWR VGND clk _01031_ reset_n keymem.key_mem\[8\]\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15271_ VGND VPWR VGND VPWR _10733_ _09988_ _10665_ _10731_ _10734_ sky130_fd_sc_hd__a31o_2
XFILLER_0_48_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24469_ VGND VPWR VPWR VGND clk _00962_ reset_n keymem.key_mem\[9\]\[78\] sky130_fd_sc_hd__dfrtp_2
X_12483_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[33\] _07578_ keymem.key_mem\[1\]\[33\]
+ _07855_ _08053_ sky130_fd_sc_hd__a22o_2
XFILLER_0_163_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17010_ VGND VPWR VGND VPWR _02758_ _02757_ _03135_ _03134_ sky130_fd_sc_hd__a21oi_2
X_14222_ _09190_ _09693_ _09060_ _09062_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_123_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_22_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14153_ VGND VPWR VGND VPWR _09623_ _09357_ _09624_ _09582_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_22_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_123_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13104_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[93\] _08577_ _08613_ _08609_ _08614_
+ sky130_fd_sc_hd__o22a_2
X_14084_ VGND VPWR VGND VPWR _09450_ _09302_ _09555_ _09397_ sky130_fd_sc_hd__a21oi_2
X_18961_ VPWR VGND _04796_ _04795_ enc_block.round_key\[53\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_21_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_123_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13035_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[87\] _07649_ keymem.key_mem\[14\]\[87\]
+ _07685_ _08551_ sky130_fd_sc_hd__a22o_2
X_17912_ VGND VPWR VGND VPWR _03872_ _03675_ _03792_ key[223] sky130_fd_sc_hd__o21a_2
X_18892_ VPWR VGND _04734_ _04733_ enc_block.round_key\[46\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_197_1446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_266_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17843_ VGND VPWR VPWR VGND _03812_ key[201] keymem.prev_key1_reg\[73\] _03825_ sky130_fd_sc_hd__mux2_2
XFILLER_0_94_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17774_ VGND VPWR _00191_ _03778_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14986_ VPWR VGND VGND VPWR _10441_ _10446_ _10450_ _10437_ _10449_ sky130_fd_sc_hd__o22ai_2
X_19513_ VGND VPWR _00552_ _05156_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16725_ VGND VPWR VGND VPWR _09714_ _09713_ _10386_ _02876_ sky130_fd_sc_hd__a21o_2
X_13937_ VPWR VGND VPWR VGND _09307_ _09291_ _09321_ _09275_ _09409_ sky130_fd_sc_hd__or4_2
X_19444_ VGND VPWR VGND VPWR _05119_ keymem.key_mem_we _02480_ _05109_ _00520_ sky130_fd_sc_hd__a31o_2
X_13868_ VPWR VGND VPWR VGND _09328_ _09291_ _09339_ _09338_ _09340_ sky130_fd_sc_hd__or4_2
X_16656_ VGND VPWR VGND VPWR _02811_ _11151_ key[157] _02798_ _02810_ sky130_fd_sc_hd__a211o_2
XFILLER_0_134_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15607_ VPWR VGND VPWR VGND _11058_ _11064_ _11062_ _10780_ _11065_ sky130_fd_sc_hd__or4_2
X_12819_ VGND VPWR VGND VPWR _08357_ _08050_ keymem.key_mem\[7\]\[65\] _08354_ _08356_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_9_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_70_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19375_ VGND VPWR VPWR VGND _05067_ _05077_ keymem.key_mem\[13\]\[121\] _05078_ sky130_fd_sc_hd__mux2_2
XFILLER_0_31_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13799_ enc_block.sword_ctr_reg\[1\] _09271_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[31\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_16587_ VGND VPWR _00038_ _02744_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_169_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18326_ VPWR VGND _04225_ enc_block.block_w1_reg\[22\] enc_block.block_w3_reg\[7\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_226_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15538_ VPWR VGND VGND VPWR _10473_ _10465_ _10559_ _10997_ sky130_fd_sc_hd__nor3_2
XFILLER_0_151_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_249_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_173_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_56_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15469_ VPWR VGND VPWR VGND _10674_ _10698_ _10928_ _10927_ _10929_ sky130_fd_sc_hd__or4_2
X_18257_ VGND VPWR _04162_ _04088_ _04161_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_245_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_702 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17208_ VPWR VGND VPWR VGND _03313_ _03312_ _03310_ _02497_ _03309_ _03314_ sky130_fd_sc_hd__a221o_2
X_18188_ VPWR VGND _04099_ enc_block.block_w2_reg\[15\] enc_block.block_w2_reg\[10\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_25_584 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_212 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17139_ VGND VPWR _03252_ _03251_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_13_768 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_163_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1228 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_106_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20150_ VGND VPWR VPWR VGND _05493_ _03460_ keymem.key_mem\[10\]\[95\] _05495_ sky130_fd_sc_hd__mux2_2
XFILLER_0_141_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_947 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_100_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1008 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20081_ VGND VPWR VPWR VGND _05457_ _03173_ keymem.key_mem\[10\]\[62\] _05459_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_146_2_Right_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_239_1229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_176_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_682 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_256_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23840_ VGND VPWR VPWR VGND clk _00333_ reset_n enc_block.block_w1_reg\[25\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_217_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_58_1037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_256_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1418 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_252_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_696 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_217_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23771_ keymem.prev_key0_reg\[127\] clk _00268_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20983_ VGND VPWR VPWR VGND _05934_ _05033_ keymem.key_mem\[7\]\[100\] _05939_ sky130_fd_sc_hd__mux2_2
X_25510_ VGND VPWR VPWR VGND clk _02003_ reset_n keymem.key_mem\[1\]\[95\] sky130_fd_sc_hd__dfrtp_2
X_22722_ VGND VPWR VPWR VGND _06822_ keymem.key_mem\[0\]\[56\] _03109_ _06826_ sky130_fd_sc_hd__mux2_2
XFILLER_0_39_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_113_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25441_ VGND VPWR VPWR VGND clk _01934_ reset_n keymem.key_mem\[1\]\[26\] sky130_fd_sc_hd__dfrtp_2
X_22653_ VGND VPWR _02051_ _06797_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_113_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21604_ VGND VPWR VPWR VGND _06263_ _10369_ keymem.key_mem\[4\]\[7\] _06269_ sky130_fd_sc_hd__mux2_2
X_25372_ VGND VPWR VPWR VGND clk _01865_ reset_n keymem.key_mem\[2\]\[85\] sky130_fd_sc_hd__dfrtp_2
X_22584_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[98\] _06767_ _06766_ _05029_ _02006_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_36_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_35_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24323_ VGND VPWR VPWR VGND clk _00816_ reset_n keymem.key_mem\[10\]\[60\] sky130_fd_sc_hd__dfrtp_2
X_21535_ VGND VPWR _06231_ _06115_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_8_784 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_860 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_62_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_562 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24254_ VGND VPWR VPWR VGND clk _00747_ reset_n keymem.key_mem\[11\]\[119\] sky130_fd_sc_hd__dfrtp_2
X_21466_ VGND VPWR VPWR VGND _06184_ _03251_ keymem.key_mem\[5\]\[71\] _06195_ sky130_fd_sc_hd__mux2_2
XFILLER_0_224_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23205_ VGND VPWR _07095_ _07092_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20417_ VGND VPWR _00976_ _05636_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24185_ VGND VPWR VPWR VGND clk _00678_ reset_n keymem.key_mem\[11\]\[50\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_181_1269 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_160_386 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21397_ VGND VPWR VPWR VGND _06151_ _02934_ keymem.key_mem\[5\]\[38\] _06159_ sky130_fd_sc_hd__mux2_2
X_23136_ VGND VPWR _02282_ _07049_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20348_ VGND VPWR _00943_ _05600_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_247_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_969 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_259_295 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_120_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23067_ VGND VPWR _02255_ _07007_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_257_1307 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20279_ VGND VPWR _00910_ _05564_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22018_ VGND VPWR VPWR VGND _06462_ _04986_ keymem.key_mem\[3\]\[72\] _06490_ sky130_fd_sc_hd__mux2_2
XFILLER_0_200_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14840_ VPWR VGND VPWR VGND _10128_ _10305_ _10304_ _09581_ sky130_fd_sc_hd__or3b_2
XFILLER_0_243_696 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14771_ VPWR VGND VGND VPWR _09411_ _09452_ _09355_ _09333_ _10237_ _10236_ sky130_fd_sc_hd__o221a_2
XFILLER_0_8_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23969_ VGND VPWR VPWR VGND clk _00462_ reset_n keymem.key_mem\[13\]\[90\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_216_1037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11983_ VGND VPWR _07586_ _07585_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13722_ VGND VPWR VGND VPWR _09194_ _09040_ _09041_ _08958_ _09010_ sky130_fd_sc_hd__a211o_2
XFILLER_0_233_1340 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_230_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16510_ VGND VPWR VGND VPWR _09505_ keymem.round_ctr_reg\[0\] _02670_ _09429_ sky130_fd_sc_hd__nand3_2
X_25708_ keymem.prev_key1_reg\[24\] clk _02201_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_17490_ VGND VPWR VPWR VGND _10366_ _11441_ key[112] _03562_ sky130_fd_sc_hd__mux2_2
XFILLER_0_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13653_ VGND VPWR _09125_ _09124_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16441_ VGND VPWR VPWR VGND _02603_ _02600_ _02599_ _09523_ _02602_ sky130_fd_sc_hd__o31ai_2
X_25639_ VGND VPWR VPWR VGND clk _02132_ reset_n keymem.key_mem\[0\]\[96\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_195_261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12604_ VGND VPWR VGND VPWR _07691_ keymem.key_mem\[3\]\[44\] _08159_ _08161_ _08163_
+ _08162_ sky130_fd_sc_hd__a2111o_2
X_16372_ VPWR VGND VPWR VGND _11615_ _02534_ _02529_ _11277_ _02535_ sky130_fd_sc_hd__or4_2
XFILLER_0_54_602 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19160_ VPWR VGND keymem.key_mem_we _04941_ _02985_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13584_ VGND VPWR _09056_ _09007_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_155_158 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15323_ VGND VPWR VGND VPWR _10785_ _10776_ _10562_ _10780_ _10784_ sky130_fd_sc_hd__a211o_2
X_18111_ VPWR VGND _04029_ _04028_ enc_block.round_key\[100\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_155_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_143_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_38_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12535_ VPWR VGND VPWR VGND _08099_ keymem.key_mem\[10\]\[38\] _07909_ keymem.key_mem\[8\]\[38\]
+ _07929_ _08100_ sky130_fd_sc_hd__a221o_2
X_19091_ VPWR VGND keymem.key_mem\[13\]\[15\] _04900_ _04887_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_227_1111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_87_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_128 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15254_ VGND VPWR VGND VPWR _10611_ _10559_ _10717_ _10521_ sky130_fd_sc_hd__a21oi_2
X_18042_ VPWR VGND VGND VPWR _03964_ enc_block.block_w3_reg\[7\] _03962_ sky130_fd_sc_hd__nand2_2
X_12466_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[32\] _07579_ keymem.key_mem\[8\]\[32\]
+ _07878_ _08037_ sky130_fd_sc_hd__a22o_2
XFILLER_0_41_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14205_ VGND VPWR VGND VPWR _09053_ _09149_ _09141_ _09177_ _09105_ _09676_ sky130_fd_sc_hd__o32a_2
XFILLER_0_227_1177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15185_ VGND VPWR VGND VPWR _10649_ _10519_ _10516_ _10515_ sky130_fd_sc_hd__o21a_2
XFILLER_0_2_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12397_ VGND VPWR enc_block.round_key\[25\] _07974_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14136_ VPWR VGND VPWR VGND _09362_ _09447_ _09607_ _09425_ _09495_ sky130_fd_sc_hd__a211oi_2
X_19993_ VGND VPWR _00776_ _05412_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_239_969 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18944_ VGND VPWR _04780_ enc_block.block_w3_reg\[19\] enc_block.block_w3_reg\[23\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_14067_ VPWR VGND VPWR VGND keymem.round_ctr_reg\[1\] _09539_ _09538_ keymem.round_ctr_reg\[0\]
+ sky130_fd_sc_hd__or3b_2
XFILLER_0_24_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_619 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13018_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[85\] _07610_ keymem.key_mem\[6\]\[85\]
+ _07818_ _08536_ sky130_fd_sc_hd__a22o_2
X_18875_ VGND VPWR _04718_ enc_block.block_w0_reg\[12\] _04646_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_218_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_197_1298 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_176_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17826_ VGND VPWR VPWR VGND _03812_ key[196] keymem.prev_key1_reg\[68\] _03813_ sky130_fd_sc_hd__mux2_2
XFILLER_0_98_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_2_Right_142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_206_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17757_ VGND VPWR VPWR VGND _03763_ _03768_ keymem.prev_key0_reg\[43\] _03769_ sky130_fd_sc_hd__mux2_2
X_14969_ VGND VPWR VGND VPWR enc_block.block_w2_reg\[15\] _08945_ _09022_ _10431_
+ _10433_ _10432_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_233_195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_222_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16708_ VPWR VGND VPWR VGND _02860_ _02677_ _02851_ key[159] _02723_ _02861_ sky130_fd_sc_hd__a221o_2
X_17688_ VGND VPWR VPWR VGND _03703_ _02483_ keymem.prev_key0_reg\[21\] _03722_ sky130_fd_sc_hd__mux2_2
XFILLER_0_193_209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19427_ VGND VPWR VGND VPWR _05110_ keymem.key_mem_we _10977_ _05109_ _00512_ sky130_fd_sc_hd__a31o_2
X_16639_ VGND VPWR _02794_ keymem.prev_key0_reg\[61\] keymem.prev_key0_reg\[93\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_169_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_130_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19358_ VPWR VGND keymem.key_mem_we _05066_ _03592_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_29_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18309_ VPWR VGND _04210_ _04209_ enc_block.round_key\[117\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_210_1181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_169_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19289_ VPWR VGND keymem.key_mem\[13\]\[93\] _05020_ _04879_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_161_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21320_ VGND VPWR VPWR VGND _06117_ _09724_ keymem.key_mem\[5\]\[1\] _06119_ sky130_fd_sc_hd__mux2_2
XFILLER_0_44_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_66_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_264 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_543 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21251_ VGND VPWR VPWR VGND _06076_ _03480_ keymem.key_mem\[6\]\[98\] _06081_ sky130_fd_sc_hd__mux2_2
X_20202_ VGND VPWR VPWR VGND _05515_ _03620_ keymem.key_mem\[10\]\[120\] _05522_ sky130_fd_sc_hd__mux2_2
X_21182_ VGND VPWR VPWR VGND _06040_ _03202_ keymem.key_mem\[6\]\[65\] _06045_ sky130_fd_sc_hd__mux2_2
XFILLER_0_106_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20133_ VGND VPWR VPWR VGND _05482_ _03393_ keymem.key_mem\[10\]\[87\] _05486_ sky130_fd_sc_hd__mux2_2
XFILLER_0_106_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20064_ VGND VPWR VPWR VGND _05446_ _03091_ keymem.key_mem\[10\]\[54\] _05450_ sky130_fd_sc_hd__mux2_2
X_24941_ VGND VPWR VPWR VGND clk _01434_ reset_n keymem.key_mem\[5\]\[38\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_147_2_Right_219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_237_490 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24872_ VGND VPWR VPWR VGND clk _01365_ reset_n keymem.key_mem\[6\]\[97\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_256_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23823_ VGND VPWR VPWR VGND clk _00316_ reset_n enc_block.block_w1_reg\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_197_548 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_75_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23754_ keymem.prev_key0_reg\[110\] clk _00251_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20966_ VPWR VGND keymem.key_mem\[7\]\[92\] _05930_ _05823_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_36_1165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22705_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[44\] _06820_ _06819_ _04943_ _02080_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_117_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23685_ keymem.prev_key0_reg\[41\] clk _00182_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20897_ VPWR VGND keymem.key_mem\[7\]\[59\] _05894_ _05886_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_222_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_187_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25424_ VGND VPWR VPWR VGND clk _01917_ reset_n keymem.key_mem\[1\]\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_996 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22636_ VGND VPWR _06789_ _03864_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_187_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_657 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_75_292 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25355_ VGND VPWR VPWR VGND clk _01848_ reset_n keymem.key_mem\[2\]\[68\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_36_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_977 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22567_ VGND VPWR VPWR VGND _06701_ keymem.key_mem\[1\]\[87\] _03393_ _06768_ sky130_fd_sc_hd__mux2_2
XFILLER_0_35_156 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_88_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_63_476 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24306_ VGND VPWR VPWR VGND clk _00799_ reset_n keymem.key_mem\[10\]\[43\] sky130_fd_sc_hd__dfrtp_2
X_12320_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[19\] _07843_ keymem.key_mem\[8\]\[19\]
+ _07903_ _07904_ sky130_fd_sc_hd__a22o_2
XFILLER_0_49_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21518_ VGND VPWR _01491_ _06222_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_228_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25286_ VGND VPWR VPWR VGND clk _01779_ reset_n keymem.key_mem\[3\]\[127\] sky130_fd_sc_hd__dfrtp_2
X_22498_ VGND VPWR _01955_ _06738_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_50_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24237_ VGND VPWR VPWR VGND clk _00730_ reset_n keymem.key_mem\[11\]\[102\] sky130_fd_sc_hd__dfrtp_2
X_12251_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[14\] _07721_ keymem.key_mem\[6\]\[14\]
+ _07712_ _07840_ sky130_fd_sc_hd__a22o_2
X_21449_ VGND VPWR _01458_ _06186_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_228_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1164 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24168_ VGND VPWR VPWR VGND clk _00661_ reset_n keymem.key_mem\[11\]\[33\] sky130_fd_sc_hd__dfrtp_2
X_12182_ VGND VPWR enc_block.round_key\[9\] _07775_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_124_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23119_ VGND VPWR VGND VPWR _02276_ _07038_ _07010_ keymem.prev_key1_reg\[99\] sky130_fd_sc_hd__o21a_2
XFILLER_0_21_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_1_Left_368 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24099_ VGND VPWR VPWR VGND clk _00592_ reset_n keymem.key_mem\[12\]\[92\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_198_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16990_ VPWR VGND VPWR VGND _03117_ _10086_ _03114_ _03115_ _03116_ _10096_ sky130_fd_sc_hd__o311a_2
XFILLER_0_159_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_101_294 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_263_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15941_ VPWR VGND VGND VPWR _11397_ _11224_ _11396_ sky130_fd_sc_hd__nand2_2
XFILLER_0_159_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18660_ _04523_ _04525_ _04294_ _04524_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_95_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15872_ VPWR VGND VPWR VGND _11206_ _11208_ _11207_ _11225_ _11328_ sky130_fd_sc_hd__or4_2
XFILLER_0_235_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17611_ VPWR VGND VPWR VGND _03667_ _03664_ _03663_ key[255] _08929_ _03668_ sky130_fd_sc_hd__a221o_2
X_14823_ VGND VPWR VGND VPWR _09749_ _09388_ _09576_ _10288_ sky130_fd_sc_hd__a21o_2
X_18591_ VPWR VGND VPWR VGND _04463_ _04401_ _04462_ sky130_fd_sc_hd__or2_2
XFILLER_0_235_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17542_ VGND VPWR VPWR VGND _03593_ keymem.key_mem\[14\]\[118\] _03607_ _03608_ sky130_fd_sc_hd__mux2_2
X_14754_ VGND VPWR VGND VPWR _09156_ _09069_ _09050_ _09203_ _10220_ sky130_fd_sc_hd__o22a_2
X_11966_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[0\] _07568_ keymem.key_mem\[6\]\[0\]
+ _07565_ _07569_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_163_1_Left_430 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_153_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13705_ VPWR VGND VGND VPWR _09177_ _08958_ _09058_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_131_2_Left_602 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14685_ VGND VPWR VGND VPWR _09204_ _09033_ _10152_ _09122_ sky130_fd_sc_hd__a21oi_2
X_17473_ VGND VPWR VPWR VGND _10378_ _03547_ key[237] _03548_ sky130_fd_sc_hd__mux2_2
X_11897_ VGND VPWR result[115] _07512_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_233_1192 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19212_ VPWR VGND keymem.key_mem\[13\]\[63\] _04973_ _04961_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16424_ VGND VPWR VGND VPWR _02573_ _02585_ _02586_ _11300_ _02575_ sky130_fd_sc_hd__nor4_2
XFILLER_0_32_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13636_ VGND VPWR _09108_ _09011_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_27_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_1085 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19143_ VPWR VGND keymem.key_mem\[13\]\[37\] _04930_ _04915_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_166_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16355_ VGND VPWR VGND VPWR _11302_ _11465_ _11351_ _11361_ _02518_ sky130_fd_sc_hd__o22a_2
XFILLER_0_54_443 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13567_ VGND VPWR _09039_ _09027_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_109_361 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_229_1228 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15306_ VPWR VGND VGND VPWR _10767_ _10768_ _10760_ sky130_fd_sc_hd__nor2_2
X_12518_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[36\] _07536_ _08084_ _08080_ _08085_
+ sky130_fd_sc_hd__o22a_2
X_16286_ VPWR VGND VGND VPWR _11303_ _02450_ _11295_ sky130_fd_sc_hd__nor2_2
X_19074_ VGND VPWR _00379_ _04890_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13498_ VGND VPWR VGND VPWR _08970_ _08968_ _08967_ keymem.prev_key1_reg\[1\] _08969_
+ _08964_ sky130_fd_sc_hd__a32o_2
XFILLER_0_246_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1406 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18025_ VPWR VGND VGND VPWR enc_block.enc_ctrl_reg\[2\] enc_block.sword_ctr_inc _07381_
+ _03947_ sky130_fd_sc_hd__nor3_2
XFILLER_0_207_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15237_ VGND VPWR VPWR VGND _10698_ _10699_ _10697_ _10700_ sky130_fd_sc_hd__or3_2
X_12449_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[30\] _07619_ keymem.key_mem\[9\]\[30\]
+ _07672_ _08022_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_244_Right_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_164_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_768 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15168_ VGND VPWR VPWR VGND _10626_ _10631_ _10621_ _10632_ sky130_fd_sc_hd__or3_2
X_14119_ VPWR VGND VGND VPWR _09480_ _09441_ _09590_ _09565_ _09404_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_227_906 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15099_ VGND VPWR _10563_ _10467_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_61_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19976_ VGND VPWR VPWR VGND _05400_ _10977_ keymem.key_mem\[10\]\[12\] _05404_ sky130_fd_sc_hd__mux2_2
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18927_ VGND VPWR _04765_ _04763_ _04764_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_126_2_Left_597 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18858_ VPWR VGND VPWR VGND _04703_ _04627_ _04702_ sky130_fd_sc_hd__or2_2
XFILLER_0_241_408 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_59_1143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_600 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_253_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1360 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17809_ VPWR VGND VGND VPWR _03801_ _03802_ _03729_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_95_1_Left_362 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18789_ VPWR VGND VPWR VGND _04641_ _04635_ _04639_ sky130_fd_sc_hd__or2_2
XFILLER_0_55_1018 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_71_2_Right_143 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20820_ VGND VPWR VGND VPWR _05852_ keymem.key_mem_we _02661_ _05850_ _01163_ sky130_fd_sc_hd__a31o_2
XFILLER_0_89_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_171_1246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_132_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20751_ VGND VPWR _01134_ _05812_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_159_261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_72_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23470_ VGND VPWR VGND VPWR _07333_ _04149_ _07093_ _07334_ enc_block.block_w3_reg\[27\]
+ sky130_fd_sc_hd__o2bb2a_2
X_20682_ VGND VPWR _01101_ _05776_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_174_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22421_ VGND VPWR VPWR VGND _06702_ keymem.key_mem\[1\]\[5\] _10194_ _06704_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_657 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25140_ VGND VPWR VPWR VGND clk _01633_ reset_n keymem.key_mem\[4\]\[109\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_936 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22352_ VGND VPWR _01881_ _06666_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_5_551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21303_ VGND VPWR VPWR VGND _06098_ _03640_ keymem.key_mem\[6\]\[123\] _06108_ sky130_fd_sc_hd__mux2_2
X_25071_ VGND VPWR VPWR VGND clk _01564_ reset_n keymem.key_mem\[4\]\[40\] sky130_fd_sc_hd__dfrtp_2
X_22283_ VGND VPWR _06630_ _03227_ _01848_ _06567_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_24022_ VGND VPWR VPWR VGND clk _00515_ reset_n keymem.key_mem\[12\]\[15\] sky130_fd_sc_hd__dfrtp_2
X_21234_ VGND VPWR VPWR VGND _06065_ _03417_ keymem.key_mem\[6\]\[90\] _06072_ sky130_fd_sc_hd__mux2_2
XFILLER_0_143_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21165_ VGND VPWR VPWR VGND _06029_ _03118_ keymem.key_mem\[6\]\[57\] _06036_ sky130_fd_sc_hd__mux2_2
XFILLER_0_223_1394 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20116_ VGND VPWR VPWR VGND _05469_ _03322_ keymem.key_mem\[10\]\[79\] _05477_ sky130_fd_sc_hd__mux2_2
X_21096_ VGND VPWR VPWR VGND _05996_ _02688_ keymem.key_mem\[6\]\[24\] _06000_ sky130_fd_sc_hd__mux2_2
XFILLER_0_217_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20047_ VGND VPWR VPWR VGND _05435_ _03015_ keymem.key_mem\[10\]\[46\] _05441_ sky130_fd_sc_hd__mux2_2
X_24924_ VGND VPWR VPWR VGND clk _01417_ reset_n keymem.key_mem\[5\]\[21\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_13_Left_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_77_1243 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_38_1205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_198_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24855_ VGND VPWR VPWR VGND clk _01348_ reset_n keymem.key_mem\[6\]\[80\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_193_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_241_953 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11820_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[13\] dec_new_block\[77\]
+ _07474_ sky130_fd_sc_hd__mux2_2
X_23806_ VGND VPWR VPWR VGND clk _00299_ reset_n enc_block.block_w0_reg\[25\] sky130_fd_sc_hd__dfrtp_2
X_24786_ VGND VPWR VPWR VGND clk _01279_ reset_n keymem.key_mem\[6\]\[11\] sky130_fd_sc_hd__dfrtp_2
X_21998_ VGND VPWR VGND VPWR _06479_ keymem.key_mem_we _03173_ _06475_ _01714_ sky130_fd_sc_hd__a31o_2
XFILLER_0_200_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_90_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_240_485 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_212_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_230_1310 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_154_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11751_ VGND VPWR result[42] _07439_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23737_ keymem.prev_key0_reg\[93\] clk _00234_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20949_ VGND VPWR VGND VPWR _05921_ keymem.key_mem_we _03356_ _05916_ _01223_ sky130_fd_sc_hd__a31o_2
XFILLER_0_230_1332 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14470_ VPWR VGND VPWR VGND _09936_ _09938_ _09937_ _09935_ _09939_ sky130_fd_sc_hd__or4_2
XFILLER_0_3_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11682_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[8\] dec_new_block\[8\]
+ _07405_ sky130_fd_sc_hd__mux2_2
X_23668_ keymem.prev_key0_reg\[24\] clk _00165_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_36_410 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_48_270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13421_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[125\] _07702_ keymem.key_mem\[11\]\[125\]
+ _07861_ _08899_ sky130_fd_sc_hd__a22o_2
XFILLER_0_165_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22619_ VGND VPWR _06779_ _06778_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25407_ VGND VPWR VPWR VGND clk _01900_ reset_n keymem.key_mem\[2\]\[120\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_49_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23599_ VGND VPWR VPWR VGND clk _00100_ reset_n keymem.key_mem\[14\]\[88\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_165_297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16140_ VPWR VGND VPWR VGND _11591_ _11593_ _11592_ _11590_ _11594_ sky130_fd_sc_hd__or4_2
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_320 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_487 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25338_ VGND VPWR VPWR VGND clk _01831_ reset_n keymem.key_mem\[2\]\[51\] sky130_fd_sc_hd__dfrtp_2
X_13352_ VPWR VGND VPWR VGND _08836_ keymem.key_mem\[13\]\[118\] _07695_ keymem.key_mem\[8\]\[118\]
+ _07958_ _08837_ sky130_fd_sc_hd__a221o_2
XFILLER_0_63_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_958 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12303_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[18\] _07622_ keymem.key_mem\[12\]\[18\]
+ _07621_ _07888_ sky130_fd_sc_hd__a22o_2
X_16071_ VPWR VGND VPWR VGND _11523_ _11525_ _11526_ _11521_ _11522_ sky130_fd_sc_hd__or4b_2
X_13283_ VPWR VGND VPWR VGND _08774_ keymem.key_mem\[11\]\[111\] _08090_ keymem.key_mem\[4\]\[111\]
+ _08077_ _08775_ sky130_fd_sc_hd__a221o_2
X_25269_ VGND VPWR VPWR VGND clk _01762_ reset_n keymem.key_mem\[3\]\[110\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_1389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_161_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15022_ VPWR VGND VGND VPWR _10480_ _10482_ _10486_ _10485_ _10484_ sky130_fd_sc_hd__o22ai_2
X_12234_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[13\] _07567_ keymem.key_mem\[10\]\[13\]
+ _07559_ _07824_ sky130_fd_sc_hd__a22o_2
XFILLER_0_32_682 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_161_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19830_ VGND VPWR VPWR VGND _05314_ keymem.key_mem\[11\]\[73\] _03268_ _05325_ sky130_fd_sc_hd__mux2_2
X_12165_ VGND VPWR _07760_ _07759_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_258_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_899 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19761_ VGND VPWR VPWR VGND _05281_ keymem.key_mem\[11\]\[40\] _02955_ _05289_ sky130_fd_sc_hd__mux2_2
XFILLER_0_159_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12096_ VGND VPWR _07694_ _07586_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16973_ VPWR VGND _03101_ _02673_ _02672_ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_198_1382 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_263_555 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18712_ VPWR VGND VPWR VGND _04571_ _04355_ _04569_ sky130_fd_sc_hd__or2_2
X_15924_ VGND VPWR _11380_ _11267_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19692_ VGND VPWR VPWR VGND _05247_ keymem.key_mem\[11\]\[7\] _10369_ _05253_ sky130_fd_sc_hd__mux2_2
X_18643_ VGND VPWR VGND VPWR _03959_ block[85] _04510_ _04509_ sky130_fd_sc_hd__a21oi_2
X_15855_ VGND VPWR _11311_ _11259_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14806_ VGND VPWR _10272_ keymem.prev_key1_reg\[6\] keymem.prev_key1_reg\[38\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_172_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18574_ _04446_ _04448_ _04065_ _04447_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_15786_ VPWR VGND VGND VPWR _11236_ _11239_ _11242_ _11211_ _11241_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_231_474 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12998_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[83\] _07597_ keymem.key_mem\[1\]\[83\]
+ _07969_ _08518_ sky130_fd_sc_hd__a22o_2
X_17525_ VGND VPWR _03593_ _09540_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14737_ VGND VPWR VGND VPWR _09211_ _09146_ _09687_ _09109_ _10203_ sky130_fd_sc_hd__o22a_2
X_11949_ VGND VPWR _07552_ _07551_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_15_1057 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17456_ VGND VPWR _03534_ _09540_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_139_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14668_ VGND VPWR VGND VPWR _09323_ _09388_ _09408_ _09466_ _10135_ sky130_fd_sc_hd__o22a_2
XFILLER_0_46_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16407_ VGND VPWR VGND VPWR _11219_ _11375_ _11460_ _11482_ _02569_ sky130_fd_sc_hd__o22a_2
XFILLER_0_116_106 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13619_ VGND VPWR _09091_ _08972_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17387_ VGND VPWR VGND VPWR _03152_ key[225] _03473_ _03474_ sky130_fd_sc_hd__a21o_2
XFILLER_0_89_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14599_ VPWR VGND VGND VPWR _09443_ _09449_ _10067_ _09380_ _09623_ sky130_fd_sc_hd__o22ai_2
X_19126_ VPWR VGND keymem.key_mem\[13\]\[31\] _04919_ _04915_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_15_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16338_ VPWR VGND VGND VPWR _11361_ _02501_ _11330_ sky130_fd_sc_hd__nor2_2
XFILLER_0_67_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19057_ VPWR VGND keymem.key_mem\[13\]\[0\] _04881_ _04880_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16269_ VGND VPWR VGND VPWR _11241_ _11344_ _11313_ _11399_ _02433_ sky130_fd_sc_hd__o22a_2
XFILLER_0_28_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_468 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_30_619 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_811 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18008_ VGND VPWR VGND VPWR _02647_ keymem.prev_key1_reg\[126\] _03679_ _03937_ sky130_fd_sc_hd__a21o_2
XFILLER_0_51_991 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_10_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19959_ VGND VPWR _00760_ _05394_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_184_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22970_ VGND VPWR VPWR VGND _02216_ _02939_ _02944_ _06925_ _06949_ sky130_fd_sc_hd__o31a_2
XFILLER_0_78_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21921_ VPWR VGND keymem.key_mem\[3\]\[27\] _06438_ _06427_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_218_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24640_ VGND VPWR VPWR VGND clk _01133_ reset_n keymem.key_mem\[8\]\[121\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_117_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21852_ VGND VPWR _01649_ _06398_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_72_2_Right_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20803_ VPWR VGND keymem.key_mem\[7\]\[16\] _05843_ _05830_ VPWR VGND sky130_fd_sc_hd__and2_2
X_24571_ VGND VPWR VPWR VGND clk _01064_ reset_n keymem.key_mem\[8\]\[52\] sky130_fd_sc_hd__dfrtp_2
X_21783_ VGND VPWR _01616_ _06362_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_77_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23522_ VGND VPWR VPWR VGND clk _00023_ reset_n keymem.key_mem\[14\]\[11\] sky130_fd_sc_hd__dfrtp_2
X_20734_ VGND VPWR _01126_ _05803_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_9_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23453_ VPWR VGND _07318_ _07256_ enc_block.block_w0_reg\[18\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_19_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20665_ VGND VPWR _01093_ _05767_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_184_1404 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22404_ VGND VPWR _01906_ _06693_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_18_498 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23384_ VGND VPWR _07257_ enc_block.block_w1_reg\[10\] _07256_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20596_ VGND VPWR _01060_ _05731_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25123_ VGND VPWR VPWR VGND clk _01616_ reset_n keymem.key_mem\[4\]\[92\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_229_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22335_ VGND VPWR _01873_ _06657_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_225_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25054_ VGND VPWR VPWR VGND clk _01547_ reset_n keymem.key_mem\[4\]\[23\] sky130_fd_sc_hd__dfrtp_2
X_22266_ VGND VPWR _01840_ _06621_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_260_1358 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1145 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_83_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_164 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24005_ VGND VPWR VPWR VGND clk _00498_ reset_n keymem.key_mem\[13\]\[126\] sky130_fd_sc_hd__dfrtp_2
X_21217_ VGND VPWR VPWR VGND _06052_ _03346_ keymem.key_mem\[6\]\[82\] _06063_ sky130_fd_sc_hd__mux2_2
XFILLER_0_130_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22197_ VGND VPWR _01807_ _06585_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_44_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_736 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21148_ VGND VPWR VPWR VGND _06018_ _03046_ keymem.key_mem\[6\]\[49\] _06027_ sky130_fd_sc_hd__mux2_2
XFILLER_0_233_706 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13970_ VPWR VGND VPWR VGND _09307_ _09290_ _09285_ _09337_ _09442_ sky130_fd_sc_hd__or4_2
XFILLER_0_232_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21079_ VGND VPWR VPWR VGND _05983_ _11446_ keymem.key_mem\[6\]\[16\] _05991_ sky130_fd_sc_hd__mux2_2
X_12921_ VGND VPWR enc_block.round_key\[75\] _08448_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24907_ VGND VPWR VPWR VGND clk _01400_ reset_n keymem.key_mem\[5\]\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_236_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_213_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15640_ VPWR VGND VPWR VGND _11097_ _09638_ _11054_ key[142] _11043_ _11098_ sky130_fd_sc_hd__a221o_2
X_24838_ VGND VPWR VPWR VGND clk _01331_ reset_n keymem.key_mem\[6\]\[63\] sky130_fd_sc_hd__dfrtp_2
X_12852_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[69\] _07779_ keymem.key_mem\[2\]\[69\]
+ _08116_ _08386_ sky130_fd_sc_hd__a22o_2
XFILLER_0_154_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_304 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11803_ VGND VPWR result[68] _07465_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_68_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15571_ VGND VPWR VGND VPWR _10184_ _10168_ _11030_ keymem.prev_key1_reg\[109\] sky130_fd_sc_hd__a21oi_2
XFILLER_0_115_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12783_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[62\] _07748_ keymem.key_mem\[11\]\[62\]
+ _08011_ _08324_ sky130_fd_sc_hd__a22o_2
X_24769_ VGND VPWR VPWR VGND clk _01262_ reset_n keymem.key_mem\[7\]\[122\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_55_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17310_ VGND VPWR VGND VPWR _11624_ _03403_ _02696_ _02701_ _03405_ sky130_fd_sc_hd__a31o_2
X_11734_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[2\] dec_new_block\[34\]
+ _07431_ sky130_fd_sc_hd__mux2_2
XFILLER_0_90_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14522_ VPWR VGND VPWR VGND _09990_ _09638_ _09929_ key[131] _09544_ _09991_ sky130_fd_sc_hd__a221o_2
XFILLER_0_51_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18290_ VPWR VGND VPWR VGND _04192_ _04189_ _04188_ enc_block.block_w0_reg\[19\]
+ _04097_ _00293_ sky130_fd_sc_hd__a221o_2
XFILLER_0_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17241_ VGND VPWR VGND VPWR _03342_ keymem.prev_key0_reg\[82\] _09795_ _11622_ _03343_
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_193_370 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14453_ VGND VPWR VGND VPWR _09912_ _09368_ _09917_ _09919_ _09922_ _09921_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_83_368 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11665_ VGND VPWR dec_next _07396_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_138_286 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13404_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[123\] _07644_ _08883_ _08877_ _08884_
+ sky130_fd_sc_hd__o22a_2
X_14384_ _09851_ _09854_ keymem.prev_key0_reg\[98\] _09852_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_17172_ VGND VPWR _03281_ _03211_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16123_ VPWR VGND VPWR VGND _11574_ _11576_ _11577_ _11388_ _11507_ sky130_fd_sc_hd__or4b_2
XFILLER_0_106_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13335_ VGND VPWR enc_block.round_key\[116\] _08821_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_52_777 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16054_ VGND VPWR VPWR VGND _11230_ _11508_ _11509_ _11338_ _11340_ sky130_fd_sc_hd__o211a_2
X_13266_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[109\] _08124_ _08759_ _08755_ _08760_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_122_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15005_ VGND VPWR _10469_ _10468_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_126_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12217_ VGND VPWR _07808_ _07807_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_161_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13197_ VPWR VGND VPWR VGND _08696_ keymem.key_mem\[5\]\[103\] _07780_ keymem.key_mem\[9\]\[103\]
+ _07593_ _08697_ sky130_fd_sc_hd__a221o_2
XFILLER_0_248_360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_23_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19813_ VGND VPWR _00692_ _05316_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_62_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12148_ VGND VPWR _07744_ _07582_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_138_58 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19744_ VGND VPWR VPWR VGND _05270_ keymem.key_mem\[11\]\[32\] _02873_ _05280_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_10_Right_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16956_ VGND VPWR VGND VPWR _02592_ _02591_ _02864_ _03086_ sky130_fd_sc_hd__a21o_2
X_12079_ VGND VPWR enc_block.round_key\[3\] _07678_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_251_514 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15907_ VPWR VGND VPWR VGND _11359_ _11362_ _11363_ _11355_ _11358_ sky130_fd_sc_hd__or4b_2
X_19675_ VGND VPWR _05243_ _05242_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_154_13 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16887_ VPWR VGND VPWR VGND _03023_ _02497_ _03019_ key[175] _02723_ _03024_ sky130_fd_sc_hd__a221o_2
XFILLER_0_188_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18626_ VPWR VGND VGND VPWR _04380_ _04495_ _04191_ sky130_fd_sc_hd__nor2_2
XFILLER_0_256_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15838_ VPWR VGND VPWR VGND _11173_ _11216_ _11179_ _11233_ _11294_ sky130_fd_sc_hd__or4_2
XFILLER_0_133_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_172_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1084 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18557_ VPWR VGND VGND VPWR _04380_ _04433_ _04116_ sky130_fd_sc_hd__nor2_2
XFILLER_0_73_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15769_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[23\] _10402_ _11225_ _09255_ _11185_
+ _11186_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_133_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17508_ VGND VPWR VGND VPWR _03578_ _03577_ _03576_ _10092_ sky130_fd_sc_hd__o21a_2
XFILLER_0_34_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_398 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18488_ VPWR VGND VGND VPWR _04328_ _04371_ _04042_ sky130_fd_sc_hd__nor2_2
XFILLER_0_191_307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17439_ VGND VPWR VPWR VGND _03467_ keymem.key_mem\[14\]\[104\] _03518_ _03519_ sky130_fd_sc_hd__mux2_2
XFILLER_0_170_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_1190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20450_ VGND VPWR VPWR VGND _05649_ _03543_ keymem.key_mem\[9\]\[108\] _05654_ sky130_fd_sc_hd__mux2_2
XFILLER_0_104_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19109_ VPWR VGND keymem.key_mem\[13\]\[23\] _04910_ _04903_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_179_21 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20381_ VPWR VGND VGND VPWR _05618_ keymem.key_mem\[9\]\[75\] _05532_ sky130_fd_sc_hd__nand2_2
XFILLER_0_3_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_207_1142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22120_ VGND VPWR _01772_ _06543_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_144_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_140_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22051_ VGND VPWR VGND VPWR _06507_ keymem.key_mem_we _03393_ _06498_ _01739_ sky130_fd_sc_hd__a31o_2
XFILLER_0_144_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_242_1099 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_80_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21002_ VGND VPWR VPWR VGND _05945_ _05052_ keymem.key_mem\[7\]\[109\] _05949_ sky130_fd_sc_hd__mux2_2
X_25810_ keymem.prev_key1_reg\[126\] clk _02303_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_255_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22953_ VGND VPWR VGND VPWR _02878_ _02876_ _02882_ _06939_ sky130_fd_sc_hd__a21o_2
X_25741_ keymem.prev_key1_reg\[57\] clk _02234_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_21904_ VPWR VGND keymem.key_mem\[3\]\[19\] _06429_ _06427_ VPWR VGND sky130_fd_sc_hd__and2_2
X_22884_ VGND VPWR _02183_ _06896_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25672_ VGND VPWR VPWR VGND clk _02165_ reset_n keymem.rcon_logic.tmp_rcon\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_151_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24623_ VGND VPWR VPWR VGND clk _01116_ reset_n keymem.key_mem\[8\]\[104\] sky130_fd_sc_hd__dfrtp_2
X_21835_ VGND VPWR VPWR VGND _06388_ _03600_ keymem.key_mem\[4\]\[117\] _06390_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_73_2_Right_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_91_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_167_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_65_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24554_ VGND VPWR VPWR VGND clk _01047_ reset_n keymem.key_mem\[8\]\[35\] sky130_fd_sc_hd__dfrtp_2
X_21766_ VGND VPWR _01608_ _06353_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_52_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_231_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23505_ VGND VPWR VPWR VGND _07093_ enc_block.block_w3_reg\[31\] _07364_ _07365_
+ sky130_fd_sc_hd__mux2_2
X_20717_ VGND VPWR VPWR VGND _05794_ _03533_ keymem.key_mem\[8\]\[106\] _05795_ sky130_fd_sc_hd__mux2_2
XFILLER_0_175_370 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_110_1_Left_377 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24485_ VGND VPWR VPWR VGND clk _00978_ reset_n keymem.key_mem\[9\]\[94\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_65_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21697_ VGND VPWR _01575_ _06317_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23436_ VGND VPWR _07304_ enc_block.round_key\[23\] _07303_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20648_ VGND VPWR _01085_ _05758_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_262_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_906 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23367_ _07240_ _07242_ _04064_ _07241_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_20579_ VGND VPWR _01052_ _05722_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_416 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13120_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[95\] _07984_ keymem.key_mem\[10\]\[95\]
+ _07876_ _08628_ sky130_fd_sc_hd__a22o_2
XFILLER_0_103_131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22318_ VGND VPWR VPWR VGND _06647_ _03374_ keymem.key_mem\[2\]\[85\] _06649_ sky130_fd_sc_hd__mux2_2
X_25106_ VGND VPWR VPWR VGND clk _01599_ reset_n keymem.key_mem\[4\]\[75\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_249_124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_162_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23298_ VGND VPWR VGND VPWR _07180_ _03981_ _07179_ _07178_ sky130_fd_sc_hd__and3b_2
XFILLER_0_123_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13051_ VGND VPWR VGND VPWR _08566_ _07737_ keymem.key_mem\[1\]\[88\] _08563_ _08565_
+ sky130_fd_sc_hd__a211o_2
X_25037_ VGND VPWR VPWR VGND clk _01530_ reset_n keymem.key_mem\[4\]\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_44_1050 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22249_ VGND VPWR VPWR VGND _06611_ _03075_ keymem.key_mem\[2\]\[52\] _06613_ sky130_fd_sc_hd__mux2_2
XFILLER_0_239_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_994 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12002_ VPWR VGND VPWR VGND _07604_ keymem.key_mem\[5\]\[0\] _07597_ keymem.key_mem\[9\]\[0\]
+ _07593_ _07605_ sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_140_2_Left_611 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_245_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_218_566 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16810_ VPWR VGND VGND VPWR _02954_ key[168] _10838_ sky130_fd_sc_hd__nand2_2
X_17790_ VGND VPWR _03788_ _03729_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_396 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16741_ VPWR VGND VPWR VGND _09855_ _02891_ _09858_ _11624_ sky130_fd_sc_hd__or3b_2
X_13953_ VPWR VGND VGND VPWR _09425_ _09303_ _09299_ sky130_fd_sc_hd__nand2_2
XFILLER_0_195_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19460_ VGND VPWR _05128_ _05094_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12904_ VPWR VGND VPWR VGND _08432_ keymem.key_mem\[13\]\[74\] _07622_ keymem.key_mem\[4\]\[74\]
+ _07914_ _08433_ sky130_fd_sc_hd__a221o_2
XFILLER_0_199_974 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16672_ VGND VPWR _02826_ _02823_ _02825_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_13884_ VPWR VGND VPWR VGND _09261_ _09317_ _09266_ _09296_ _09356_ sky130_fd_sc_hd__or4_2
X_18411_ VPWR VGND VGND VPWR _04301_ _04302_ _03974_ sky130_fd_sc_hd__nor2_2
X_15623_ VPWR VGND VGND VPWR _10761_ _10762_ _10766_ _11081_ sky130_fd_sc_hd__nor3_2
X_12835_ VGND VPWR VGND VPWR _07610_ keymem.key_mem\[7\]\[67\] _08368_ _08370_ _08371_
+ _07662_ sky130_fd_sc_hd__a2111o_2
X_19391_ VGND VPWR _00498_ _05088_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_29_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_1141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_1190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18342_ VGND VPWR VGND VPWR _09505_ _09429_ _04073_ _04240_ sky130_fd_sc_hd__a21o_2
X_15554_ VGND VPWR VGND VPWR _10476_ _10490_ _10459_ _10477_ _10514_ _11013_ sky130_fd_sc_hd__o32a_2
XFILLER_0_33_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12766_ VGND VPWR VGND VPWR _07778_ keymem.key_mem\[3\]\[60\] _08306_ _08308_ _08309_
+ _08243_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_12_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_189_1145 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_204_Right_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14505_ VGND VPWR VGND VPWR _09154_ _09148_ _08999_ _09105_ _09071_ _09974_ sky130_fd_sc_hd__o32a_2
X_11717_ VGND VPWR result[25] _07422_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18273_ VPWR VGND VPWR VGND _04176_ block[114] _04076_ enc_block.block_w1_reg\[18\]
+ _04171_ _04177_ sky130_fd_sc_hd__a221o_2
X_15485_ VGND VPWR VGND VPWR _10867_ _10944_ _10635_ _10945_ sky130_fd_sc_hd__a21o_2
X_12697_ VPWR VGND VPWR VGND _08246_ keymem.key_mem\[7\]\[53\] _07703_ keymem.key_mem\[10\]\[53\]
+ _07743_ _08247_ sky130_fd_sc_hd__a221o_2
XFILLER_0_12_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_210_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_140_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_722 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17224_ VPWR VGND VPWR VGND _03327_ _03325_ _10096_ _03324_ _03328_ sky130_fd_sc_hd__a22o_2
X_14436_ VGND VPWR VGND VPWR _09380_ _09440_ _09475_ _09495_ _09905_ sky130_fd_sc_hd__o22a_2
X_11648_ VPWR VGND VPWR VGND _07385_ keymem.round_ctr_reg\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_71_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17155_ VPWR VGND VPWR VGND _03265_ _03262_ _09534_ _03261_ _03266_ sky130_fd_sc_hd__a22o_2
X_14367_ VGND VPWR VGND VPWR _09160_ _09109_ _09224_ _09837_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_141_248 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16106_ VPWR VGND _11560_ keymem.prev_key0_reg\[82\] keymem.prev_key0_reg\[50\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
X_13318_ VPWR VGND VPWR VGND _08805_ keymem.key_mem\[14\]\[115\] _08032_ keymem.key_mem\[4\]\[115\]
+ _07637_ _08806_ sky130_fd_sc_hd__a221o_2
X_14298_ VPWR VGND VPWR VGND _09767_ _09768_ _09765_ _09766_ sky130_fd_sc_hd__or3b_2
X_17086_ VGND VPWR VPWR VGND _09732_ _09792_ key[194] _03204_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_72_2_Left_543 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_204_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16037_ VGND VPWR VGND VPWR _11492_ _11434_ _11409_ _11491_ _11271_ sky130_fd_sc_hd__a211o_2
XFILLER_0_23_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13249_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[108\] _07659_ keymem.key_mem\[7\]\[108\]
+ _07608_ _08744_ sky130_fd_sc_hd__a22o_2
XFILLER_0_255_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_460 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_27_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_213_Right_82 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_196_1105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_58_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17988_ VGND VPWR VPWR VGND _03674_ _03923_ keymem.prev_key0_reg\[119\] _03924_ sky130_fd_sc_hd__mux2_2
XFILLER_0_252_823 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_165_23 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_694 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_224_536 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_178_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_97_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19727_ VGND VPWR _00651_ _05271_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16939_ VGND VPWR VGND VPWR _03071_ _10328_ _02877_ key[52] sky130_fd_sc_hd__o21a_2
X_19658_ VGND VPWR VPWR VGND _05227_ _05077_ keymem.key_mem\[12\]\[121\] _05233_ sky130_fd_sc_hd__mux2_2
X_18609_ VPWR VGND _04479_ enc_block.block_w1_reg\[26\] enc_block.block_w2_reg\[17\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_172_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19589_ VGND VPWR VPWR VGND _05183_ _05013_ keymem.key_mem\[12\]\[88\] _05197_ sky130_fd_sc_hd__mux2_2
XFILLER_0_149_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_825 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_34_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_222_Right_91 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21620_ VGND VPWR _01538_ _06277_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_133_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21551_ VGND VPWR _01507_ _06239_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_379 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20502_ VGND VPWR _01015_ _05682_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24270_ VGND VPWR VPWR VGND clk _00763_ reset_n keymem.key_mem\[10\]\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_7_465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21482_ VGND VPWR _01474_ _06203_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_476 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_69_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_209_1215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_132_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23221_ VGND VPWR _07110_ _07108_ _07109_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20433_ VGND VPWR VPWR VGND _05638_ _03492_ keymem.key_mem\[9\]\[100\] _05645_ sky130_fd_sc_hd__mux2_2
XFILLER_0_43_574 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_99_95 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_200_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23152_ VGND VPWR _02287_ _07060_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20364_ VGND VPWR VPWR VGND _05602_ _03217_ keymem.key_mem\[9\]\[67\] _05609_ sky130_fd_sc_hd__mux2_2
XFILLER_0_222_1415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22103_ VGND VPWR _01764_ _06534_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23083_ VGND VPWR VGND VPWR _07017_ _03370_ _03369_ _03373_ _07011_ sky130_fd_sc_hd__a211o_2
XFILLER_0_105_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20295_ VGND VPWR VPWR VGND _05569_ _02894_ keymem.key_mem\[9\]\[34\] _05573_ sky130_fd_sc_hd__mux2_2
XFILLER_0_45_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_144_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22034_ VPWR VGND keymem.key_mem\[3\]\[79\] _06499_ _06484_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_80_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_609 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_834 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_76_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_242_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23985_ VGND VPWR VPWR VGND clk _00478_ reset_n keymem.key_mem\[13\]\[106\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_225_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25724_ keymem.prev_key1_reg\[40\] clk _02217_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22936_ VGND VPWR VGND VPWR _02732_ _06928_ _02741_ _06929_ sky130_fd_sc_hd__a21o_2
XFILLER_0_151_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25655_ VGND VPWR VPWR VGND clk _02148_ reset_n keymem.key_mem\[0\]\[112\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_155_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22867_ VGND VPWR VGND VPWR _06885_ _09636_ _03795_ _06884_ _09723_ sky130_fd_sc_hd__a211o_2
XFILLER_0_196_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_836 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_52_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24606_ VGND VPWR VPWR VGND clk _01099_ reset_n keymem.key_mem\[8\]\[87\] sky130_fd_sc_hd__dfrtp_2
X_12620_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[46\] _07592_ keymem.key_mem\[11\]\[46\]
+ _07861_ _08177_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_74_2_Right_146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21818_ VGND VPWR VPWR VGND _06377_ _03550_ keymem.key_mem\[4\]\[109\] _06381_ sky130_fd_sc_hd__mux2_2
XFILLER_0_196_999 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25586_ VGND VPWR VPWR VGND clk _02079_ reset_n keymem.key_mem\[0\]\[43\] sky130_fd_sc_hd__dfrtp_2
X_22798_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[101\] _06850_ _06849_ _05035_ _02137_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_112_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12551_ VGND VPWR enc_block.round_key\[39\] _08114_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_368 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21749_ VGND VPWR VPWR VGND _06344_ _03295_ keymem.key_mem\[4\]\[76\] _06345_ sky130_fd_sc_hd__mux2_2
X_24537_ VGND VPWR VPWR VGND clk _01030_ reset_n keymem.key_mem\[8\]\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_828 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_87_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_241_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_582 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_266_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12482_ VGND VPWR _08052_ _07724_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15270_ VPWR VGND VGND VPWR _10732_ _10733_ key[9] sky130_fd_sc_hd__nor2_2
X_24468_ VGND VPWR VPWR VGND clk _00961_ reset_n keymem.key_mem\[9\]\[77\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_46_390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_87_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14221_ VGND VPWR VGND VPWR _09691_ _09690_ _09692_ _09689_ _09688_ sky130_fd_sc_hd__nand4_2
X_23419_ VGND VPWR _07289_ enc_block.round_key\[21\] _07288_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_168 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_266_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24399_ VGND VPWR VPWR VGND clk _00892_ reset_n keymem.key_mem\[9\]\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_110_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_22_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14152_ VGND VPWR _09623_ _09622_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_85_1172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_127_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_162_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13103_ VGND VPWR VGND VPWR _08613_ _07580_ keymem.key_mem\[12\]\[93\] _08610_ _08612_
+ sky130_fd_sc_hd__a211o_2
X_14083_ _09552_ _09554_ _09370_ _09553_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_18960_ VPWR VGND VPWR VGND _04794_ block[53] _04744_ enc_block.block_w3_reg\[21\]
+ _04666_ _04795_ sky130_fd_sc_hd__a221o_2
XFILLER_0_123_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_162_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13034_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[87\] _07779_ keymem.key_mem\[6\]\[87\]
+ _07657_ _08550_ sky130_fd_sc_hd__a22o_2
X_17911_ VGND VPWR VGND VPWR _03732_ keymem.prev_key1_reg\[95\] _03864_ _03871_ sky130_fd_sc_hd__a21o_2
XPHY_EDGE_ROW_5_Left_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18891_ VPWR VGND VPWR VGND _04732_ block[46] _04351_ enc_block.block_w0_reg\[14\]
+ _03978_ _04733_ sky130_fd_sc_hd__a221o_2
XFILLER_0_123_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17842_ VGND VPWR _00213_ _03824_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_98_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_266_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_94_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17773_ VGND VPWR VPWR VGND _03777_ _03052_ keymem.prev_key0_reg\[50\] _03778_ sky130_fd_sc_hd__mux2_2
X_14985_ VGND VPWR _10449_ _10448_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_234_878 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_238_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19512_ VGND VPWR VPWR VGND _05151_ _04958_ keymem.key_mem\[12\]\[52\] _05156_ sky130_fd_sc_hd__mux2_2
X_16724_ VGND VPWR _02875_ _09543_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13936_ VGND VPWR _09408_ _09407_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_214_580 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_134_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19443_ VPWR VGND keymem.key_mem\[12\]\[20\] _05119_ _05116_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_88_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16655_ VGND VPWR VPWR VGND _02810_ _02708_ _02806_ _02807_ _02809_ sky130_fd_sc_hd__o31a_2
X_13867_ VGND VPWR _09339_ _09321_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_173_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15606_ VPWR VGND VPWR VGND _10984_ _11063_ _11064_ _10886_ _10871_ sky130_fd_sc_hd__or4b_2
XFILLER_0_134_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_324 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12818_ VPWR VGND VPWR VGND _08355_ keymem.key_mem\[5\]\[65\] _08052_ keymem.key_mem\[3\]\[65\]
+ _07690_ _08356_ sky130_fd_sc_hd__a221o_2
X_19374_ VPWR VGND keymem.key_mem_we _05077_ _03627_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_158_156 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16586_ VGND VPWR VPWR VGND _02662_ keymem.key_mem\[14\]\[26\] _02743_ _02744_ sky130_fd_sc_hd__mux2_2
X_13798_ VPWR VGND VGND VPWR enc_block.block_w1_reg\[31\] enc_block.sword_ctr_reg\[0\]
+ _09270_ sky130_fd_sc_hd__or2b_2
XFILLER_0_70_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_806 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18325_ VPWR VGND VPWR VGND _04224_ _04189_ _04222_ enc_block.block_w0_reg\[22\]
+ _04097_ _00296_ sky130_fd_sc_hd__a221o_2
XFILLER_0_169_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15537_ VPWR VGND VGND VPWR _10587_ _10996_ _10488_ sky130_fd_sc_hd__nor2_2
X_12749_ VPWR VGND VPWR VGND _08293_ keymem.key_mem\[10\]\[58\] _07876_ keymem.key_mem\[8\]\[58\]
+ _07541_ _08294_ sky130_fd_sc_hd__a221o_2
XFILLER_0_44_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_38_891 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18256_ VPWR VGND _04161_ enc_block.block_w1_reg\[23\] enc_block.block_w1_reg\[16\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_71_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15468_ VPWR VGND VGND VPWR _10628_ _10928_ _10522_ sky130_fd_sc_hd__nor2_2
X_17207_ key[206] _03313_ keylen _10967_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_14419_ VGND VPWR VGND VPWR _09410_ _09401_ _09888_ _09399_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_114_226 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_245_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18187_ VPWR VGND _04098_ _04022_ enc_block.block_w3_reg\[2\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15399_ VGND VPWR VPWR VGND _10859_ _10860_ _10857_ _10856_ _10511_ _10541_ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_13_714 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17138_ VPWR VGND VPWR VGND _03250_ _02497_ _03247_ key[199] _03211_ _03251_ sky130_fd_sc_hd__a221o_2
XFILLER_0_52_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_180_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1183 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_229_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17069_ VGND VPWR VGND VPWR _09508_ keymem.prev_key0_reg\[64\] _03189_ _08937_ sky130_fd_sc_hd__nand3_2
XFILLER_0_229_628 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_141_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_11 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20080_ VGND VPWR _00817_ _05458_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_141_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1208 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_120_1_Right_721 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_225_801 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_221_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_85_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_256_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_719 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23770_ keymem.prev_key0_reg\[126\] clk _00267_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20982_ VGND VPWR _01239_ _05938_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_189_270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22721_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[55\] _06820_ _06819_ _04963_ _02091_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_152_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_113_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25440_ VGND VPWR VPWR VGND clk _01933_ reset_n keymem.key_mem\[1\]\[25\] sky130_fd_sc_hd__dfrtp_2
X_22652_ VGND VPWR VPWR VGND _06785_ keymem.key_mem\[0\]\[15\] _11149_ _06797_ sky130_fd_sc_hd__mux2_2
XFILLER_0_152_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_250_1176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_87_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21603_ VGND VPWR _01530_ _06268_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_258_Right_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25371_ VGND VPWR VPWR VGND clk _01864_ reset_n keymem.key_mem\[2\]\[84\] sky130_fd_sc_hd__dfrtp_2
X_22583_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[97\] _06767_ _06766_ _05027_ _02005_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_1_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24322_ VGND VPWR VPWR VGND clk _00815_ reset_n keymem.key_mem\[10\]\[59\] sky130_fd_sc_hd__dfrtp_2
X_21534_ VGND VPWR _01499_ _06230_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_1_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_69_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_105_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_796 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_62_146 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24253_ VGND VPWR VPWR VGND clk _00746_ reset_n keymem.key_mem\[11\]\[118\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_7_295 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21465_ VGND VPWR _01466_ _06194_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_263_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23204_ VGND VPWR VGND VPWR _07091_ _03992_ _07094_ _02305_ sky130_fd_sc_hd__a21o_2
XFILLER_0_181_1237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_382 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20416_ VGND VPWR VPWR VGND _05627_ _03435_ keymem.key_mem\[9\]\[92\] _05636_ sky130_fd_sc_hd__mux2_2
XFILLER_0_43_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24184_ VGND VPWR VPWR VGND clk _00677_ reset_n keymem.key_mem\[11\]\[49\] sky130_fd_sc_hd__dfrtp_2
X_21396_ VGND VPWR _01433_ _06158_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23135_ VGND VPWR VPWR VGND _07032_ _07048_ keymem.prev_key1_reg\[105\] _07049_ sky130_fd_sc_hd__mux2_2
XFILLER_0_113_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20347_ VGND VPWR VPWR VGND _05591_ _03140_ keymem.key_mem\[9\]\[59\] _05600_ sky130_fd_sc_hd__mux2_2
X_23066_ VGND VPWR VPWR VGND _06992_ _07006_ keymem.prev_key1_reg\[78\] _07007_ sky130_fd_sc_hd__mux2_2
XFILLER_0_120_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20278_ VGND VPWR VPWR VGND _05558_ _02743_ keymem.key_mem\[9\]\[26\] _05564_ sky130_fd_sc_hd__mux2_2
XFILLER_0_200_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22017_ VGND VPWR VGND VPWR _06489_ keymem.key_mem_we _03252_ _06475_ _01723_ sky130_fd_sc_hd__a31o_2
XFILLER_0_215_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_200_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1043 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_242_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_255_1065 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14770_ VGND VPWR VGND VPWR _09565_ _09418_ _09349_ _09749_ _10236_ sky130_fd_sc_hd__o22a_2
X_23968_ VGND VPWR VPWR VGND clk _00461_ reset_n keymem.key_mem\[13\]\[89\] sky130_fd_sc_hd__dfrtp_2
X_11982_ VPWR VGND VGND VPWR _07554_ _07585_ _07531_ sky130_fd_sc_hd__nor2_2
XFILLER_0_59_909 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_192_1388 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13721_ VPWR VGND VPWR VGND _09193_ _09187_ _09192_ sky130_fd_sc_hd__or2_2
X_25707_ keymem.prev_key1_reg\[23\] clk _02200_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22919_ VGND VPWR VGND VPWR _02197_ _06917_ _06916_ keymem.prev_key1_reg\[20\] sky130_fd_sc_hd__o21a_2
XFILLER_0_105_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23899_ VGND VPWR VPWR VGND clk _00392_ reset_n keymem.key_mem\[13\]\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16440_ VPWR VGND VGND VPWR _02602_ keymem.prev_key1_reg\[54\] _08927_ sky130_fd_sc_hd__nand2_2
X_13652_ VGND VPWR _09124_ _09123_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25638_ VGND VPWR VPWR VGND clk _02131_ reset_n keymem.key_mem\[0\]\[95\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12603_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[44\] _07760_ keymem.key_mem\[11\]\[44\]
+ _08011_ _08162_ sky130_fd_sc_hd__a22o_2
X_16371_ VPWR VGND VPWR VGND _02531_ _02533_ _02532_ _02530_ _02534_ sky130_fd_sc_hd__or4_2
XFILLER_0_13_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_2_Right_147 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13583_ VPWR VGND VPWR VGND _09055_ _09048_ _09054_ sky130_fd_sc_hd__or2_2
X_25569_ VGND VPWR VPWR VGND clk _02062_ reset_n keymem.key_mem\[0\]\[26\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_52_1193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18110_ VPWR VGND VPWR VGND _04027_ block[100] _03959_ enc_block.block_w3_reg\[4\]
+ _03954_ _04028_ sky130_fd_sc_hd__a221o_2
X_15322_ VPWR VGND VPWR VGND _10783_ _10784_ _10781_ _10782_ sky130_fd_sc_hd__or3b_2
XFILLER_0_13_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12534_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[38\] _07716_ keymem.key_mem\[11\]\[38\]
+ _07599_ _08099_ sky130_fd_sc_hd__a22o_2
X_19090_ VGND VPWR VGND VPWR _04899_ keymem.key_mem_we _11099_ _04896_ _00386_ sky130_fd_sc_hd__a31o_2
XFILLER_0_30_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18041_ VPWR VGND VPWR VGND _03963_ enc_block.block_w3_reg\[7\] _03962_ sky130_fd_sc_hd__or2_2
XFILLER_0_87_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15253_ VPWR VGND VGND VPWR _10503_ _10524_ _10716_ _10437_ _10557_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_227_1134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_163_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12465_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[31\] _08027_ _08036_ _08031_ enc_block.round_key\[31\]
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_35_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14204_ VPWR VGND VGND VPWR _09646_ _09675_ _09200_ sky130_fd_sc_hd__nor2_2
XFILLER_0_22_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15184_ VPWR VGND VGND VPWR _10648_ _10645_ _10647_ sky130_fd_sc_hd__nand2_2
XFILLER_0_111_207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12396_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[25\] _07893_ _07973_ _07967_ _07974_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_61_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_555 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_239_926 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14135_ VGND VPWR VPWR VGND _09601_ _09605_ _09599_ _09606_ sky130_fd_sc_hd__or3_2
X_19992_ VGND VPWR VPWR VGND _05400_ _02480_ keymem.key_mem\[10\]\[20\] _05412_ sky130_fd_sc_hd__mux2_2
XFILLER_0_39_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18943_ VPWR VGND VPWR VGND _04779_ _04664_ _04777_ enc_block.block_w2_reg\[19\]
+ _04709_ _00359_ sky130_fd_sc_hd__a221o_2
X_14066_ VGND VPWR VGND VPWR keymem.round_ctr_reg\[3\] keymem.key_mem_we _09538_ keymem.round_ctr_reg\[2\]
+ sky130_fd_sc_hd__nand3_2
XFILLER_0_219_650 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13017_ VGND VPWR VGND VPWR _07842_ keymem.key_mem\[9\]\[85\] _08532_ _08534_ _08535_
+ _08020_ sky130_fd_sc_hd__a2111o_2
X_18874_ VPWR VGND VPWR VGND _04717_ _04664_ _04716_ enc_block.block_w2_reg\[12\]
+ _04709_ _00352_ sky130_fd_sc_hd__a221o_2
XFILLER_0_247_992 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_98_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_1_Left_402 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_158_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17825_ VGND VPWR _03812_ _03211_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_94_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_804 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_59_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17756_ VGND VPWR VGND VPWR _03670_ keymem.prev_key1_reg\[43\] _02982_ _03768_ sky130_fd_sc_hd__a21o_2
XFILLER_0_169_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14968_ VGND VPWR VGND VPWR _10432_ enc_block.sword_ctr_reg\[0\] enc_block.block_w1_reg\[15\]
+ enc_block.sword_ctr_reg\[1\] sky130_fd_sc_hd__and3b_2
XFILLER_0_222_848 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_178_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16707_ VPWR VGND VPWR VGND _02860_ _10325_ _02857_ _02858_ _02859_ _10281_ sky130_fd_sc_hd__o311a_2
X_13919_ VGND VPWR _09391_ _09390_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17687_ VGND VPWR _00161_ _03721_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_59_Left_327 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14899_ _10361_ _10364_ keymem.prev_key0_reg\[103\] _10362_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_19426_ VPWR VGND keymem.key_mem\[12\]\[12\] _05110_ _05102_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_9_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16638_ VPWR VGND _02793_ _02792_ keymem.prev_key0_reg\[125\] VPWR VGND sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_8_Right_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_134_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19357_ VGND VPWR _00487_ _05065_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_31_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16569_ VGND VPWR VGND VPWR _02726_ _10360_ _02724_ _02725_ _02727_ sky130_fd_sc_hd__a31o_2
XFILLER_0_17_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_485 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18308_ VPWR VGND VPWR VGND _04208_ block[117] _04076_ enc_block.block_w1_reg\[21\]
+ _04171_ _04209_ sky130_fd_sc_hd__a221o_2
X_19288_ VGND VPWR VGND VPWR _05019_ keymem.key_mem_we _03435_ _04999_ _00464_ sky130_fd_sc_hd__a31o_2
XFILLER_0_169_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18239_ VPWR VGND VPWR VGND _04145_ block[111] _04139_ enc_block.block_w2_reg\[15\]
+ _04138_ _04146_ sky130_fd_sc_hd__a221o_2
XFILLER_0_245_1223 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_111_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21250_ VGND VPWR _01365_ _06080_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_142_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20201_ VGND VPWR _00875_ _05521_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21181_ VGND VPWR _01332_ _06044_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_106_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20132_ VGND VPWR _00842_ _05485_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_39_Right_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_96_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_1_Left_334 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_238_981 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20063_ VGND VPWR _00809_ _05449_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24940_ VGND VPWR VPWR VGND clk _01433_ reset_n keymem.key_mem\[5\]\[37\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_1_Right_722 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_176_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24871_ VGND VPWR VPWR VGND clk _01364_ reset_n keymem.key_mem\[6\]\[96\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_224_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_77_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23822_ VGND VPWR VPWR VGND clk _00315_ reset_n enc_block.block_w1_reg\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_256_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_240_634 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_240_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_217_1358 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23753_ keymem.prev_key0_reg\[109\] clk _00250_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20965_ VGND VPWR VGND VPWR _05929_ keymem.key_mem_we _03427_ _05916_ _01231_ sky130_fd_sc_hd__a31o_2
XFILLER_0_67_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22704_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[43\] _06820_ _06819_ _04941_ _02079_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_36_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_238 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_48_430 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_67_249 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_113_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20896_ VGND VPWR _05893_ _05820_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23684_ keymem.prev_key0_reg\[40\] clk _00181_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_48_Right_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_49_964 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25423_ VGND VPWR VPWR VGND clk _01916_ reset_n keymem.key_mem\[1\]\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_113_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22635_ VGND VPWR _02042_ _06788_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_192_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_187_1413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_14_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_192_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22566_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[86\] _06767_ _06766_ _05010_ _01994_
+ sky130_fd_sc_hd__a22o_2
X_25354_ VGND VPWR VPWR VGND clk _01847_ reset_n keymem.key_mem\[2\]\[67\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_49_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_187_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_84_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21517_ VGND VPWR VPWR VGND _06220_ _03459_ keymem.key_mem\[5\]\[95\] _06222_ sky130_fd_sc_hd__mux2_2
XFILLER_0_267_1481 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24305_ VGND VPWR VPWR VGND clk _00798_ reset_n keymem.key_mem\[10\]\[42\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_23_308 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_179 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22497_ VGND VPWR VPWR VGND _06726_ keymem.key_mem\[1\]\[47\] _03025_ _06738_ sky130_fd_sc_hd__mux2_2
X_25285_ VGND VPWR VPWR VGND clk _01778_ reset_n keymem.key_mem\[3\]\[126\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_263_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12250_ VGND VPWR _07839_ _07838_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21448_ VGND VPWR VPWR VGND _06184_ _03172_ keymem.key_mem\[5\]\[62\] _06186_ sky130_fd_sc_hd__mux2_2
X_24236_ VGND VPWR VPWR VGND clk _00729_ reset_n keymem.key_mem\[11\]\[101\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_31_363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24167_ VGND VPWR VPWR VGND clk _00660_ reset_n keymem.key_mem\[11\]\[32\] sky130_fd_sc_hd__dfrtp_2
X_12181_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[9\] _07535_ _07774_ _07769_ _07775_
+ sky130_fd_sc_hd__o22a_2
X_21379_ VGND VPWR _01425_ _06149_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_57_Right_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23118_ VGND VPWR VGND VPWR _07038_ _03482_ _03212_ _06924_ _03484_ sky130_fd_sc_hd__a211o_2
XFILLER_0_124_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24098_ VGND VPWR VPWR VGND clk _00591_ reset_n keymem.key_mem\[12\]\[91\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_21_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15940_ VPWR VGND VGND VPWR _11396_ _11395_ _11221_ sky130_fd_sc_hd__nand2_2
X_23049_ VPWR VGND VPWR VGND _06997_ keymem.prev_key1_reg\[71\] _06926_ sky130_fd_sc_hd__or2_2
XFILLER_0_159_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_748 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15871_ VGND VPWR _11327_ _11326_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_239_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_95_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17610_ VPWR VGND VPWR VGND _03665_ _10323_ _03667_ _03666_ keylen sky130_fd_sc_hd__a211oi_2
XFILLER_0_235_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14822_ VGND VPWR _10287_ _10286_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18590_ VGND VPWR _04462_ enc_block.block_w1_reg\[24\] _04461_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17541_ VGND VPWR VGND VPWR _03152_ key[246] _03606_ _03607_ sky130_fd_sc_hd__a21o_2
XFILLER_0_235_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14753_ VGND VPWR VGND VPWR _09646_ _09159_ _09216_ _09140_ _10219_ sky130_fd_sc_hd__o22a_2
X_11965_ VGND VPWR _07568_ _07567_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_153_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13704_ VPWR VGND VGND VPWR _09176_ _09171_ _09175_ sky130_fd_sc_hd__nand2_2
X_17472_ VPWR VGND VPWR VGND _03547_ _11030_ _11031_ sky130_fd_sc_hd__or2_2
XFILLER_0_230_188 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14684_ VPWR VGND VPWR VGND _10016_ _09218_ _10149_ _10150_ _10151_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_131_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11896_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[19\] dec_new_block\[115\]
+ _07512_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_81_2_Left_552 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19211_ VGND VPWR VGND VPWR _04972_ keymem.key_mem_we _03173_ _04968_ _00434_ sky130_fd_sc_hd__a31o_2
X_16423_ VPWR VGND VPWR VGND _02579_ _02584_ _02585_ _11382_ _02578_ sky130_fd_sc_hd__or4b_2
X_13635_ VGND VPWR _09107_ _09090_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_55_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_271 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_76_2_Right_148 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19142_ VGND VPWR _00408_ _04929_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16354_ VGND VPWR VGND VPWR _02517_ _11365_ _11395_ _11390_ _11348_ _11356_ sky130_fd_sc_hd__a32o_2
XFILLER_0_41_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13566_ VPWR VGND VPWR VGND _09020_ _09037_ _09038_ _09000_ _09012_ sky130_fd_sc_hd__or4b_2
XFILLER_0_166_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_246_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15305_ VPWR VGND VPWR VGND _10762_ _10766_ _10763_ _10761_ _10767_ sky130_fd_sc_hd__or4_2
X_12517_ VGND VPWR VGND VPWR _08084_ _07721_ keymem.key_mem\[14\]\[36\] _08081_ _08083_
+ sky130_fd_sc_hd__a211o_2
X_19073_ VGND VPWR VPWR VGND _04877_ _04889_ keymem.key_mem\[13\]\[7\] _04890_ sky130_fd_sc_hd__mux2_2
X_16285_ VGND VPWR VGND VPWR _02448_ _02447_ _02449_ _02446_ _02445_ sky130_fd_sc_hd__nand4_2
XFILLER_0_26_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13497_ VGND VPWR _08969_ _08954_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_42_639 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_207_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18024_ VGND VPWR VGND VPWR _07375_ enc_block.ready _07382_ _00273_ sky130_fd_sc_hd__a21o_2
XFILLER_0_124_354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15236_ VPWR VGND VGND VPWR _10595_ _10699_ _10497_ sky130_fd_sc_hd__nor2_2
XFILLER_0_124_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_229_Left_496 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_242_1418 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12448_ VGND VPWR VGND VPWR _08016_ keymem.key_mem\[7\]\[30\] _08017_ _08019_ _08021_
+ _08020_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_23_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15167_ VGND VPWR VGND VPWR _10631_ _10574_ _10628_ _10583_ _10627_ _10630_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_22_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12379_ VGND VPWR _07958_ _07903_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_103_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14118_ VPWR VGND VGND VPWR _09557_ _09570_ _09588_ _09589_ sky130_fd_sc_hd__nor3_2
XFILLER_0_142_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15098_ VGND VPWR _10562_ _10473_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19975_ VGND VPWR _05403_ _10913_ _00767_ _05402_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_205_1295 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_103_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1030 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18926_ VGND VPWR _04764_ enc_block.block_w3_reg\[17\] enc_block.block_w2_reg\[26\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_14049_ VGND VPWR _09521_ _09510_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_238_299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_66_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_98_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18857_ VGND VPWR _04702_ _04635_ _04701_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_206_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_253_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17808_ VGND VPWR VGND VPWR _03737_ keymem.prev_key1_reg\[62\] _03801_ _03789_ sky130_fd_sc_hd__a21oi_2
X_18788_ VPWR VGND VGND VPWR _04640_ _04635_ _04639_ sky130_fd_sc_hd__nand2_2
XFILLER_0_238_1093 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_222_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_214_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17739_ VGND VPWR VPWR VGND _03723_ _03757_ keymem.prev_key0_reg\[36\] _03758_ sky130_fd_sc_hd__mux2_2
X_20750_ VGND VPWR VPWR VGND _05805_ _03633_ keymem.key_mem\[8\]\[122\] _05812_ sky130_fd_sc_hd__mux2_2
XFILLER_0_49_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_216_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19409_ VGND VPWR VGND VPWR _05100_ keymem.key_mem_we _10099_ _05093_ _00504_ sky130_fd_sc_hd__a31o_2
XFILLER_0_110_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20681_ VGND VPWR VPWR VGND _05772_ _03409_ keymem.key_mem\[8\]\[89\] _05776_ sky130_fd_sc_hd__mux2_2
XFILLER_0_58_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22420_ VGND VPWR _01912_ _06703_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_93_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22351_ VGND VPWR VPWR VGND _06658_ _03499_ keymem.key_mem\[2\]\[101\] _06666_ sky130_fd_sc_hd__mux2_2
X_21302_ VGND VPWR _01390_ _06107_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25070_ VGND VPWR VPWR VGND clk _01563_ reset_n keymem.key_mem\[4\]\[39\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_115_376 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22282_ VPWR VGND VGND VPWR _06630_ keymem.key_mem\[2\]\[68\] _06567_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1305 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_875 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_206_1037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24021_ VGND VPWR VPWR VGND clk _00514_ reset_n keymem.key_mem\[12\]\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_198_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21233_ VGND VPWR _01357_ _06071_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_223_1340 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_694 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_223_1362 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21164_ VGND VPWR _01324_ _06035_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_106_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20115_ VGND VPWR _00834_ _05476_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21095_ VGND VPWR _01291_ _05999_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20046_ VGND VPWR _00801_ _05440_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24923_ VGND VPWR VPWR VGND clk _01416_ reset_n keymem.key_mem\[5\]\[20\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_122_1_Right_723 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_99_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24854_ VGND VPWR VPWR VGND clk _01347_ reset_n keymem.key_mem\[6\]\[79\] sky130_fd_sc_hd__dfrtp_2
X_23805_ VGND VPWR VPWR VGND clk _00298_ reset_n enc_block.block_w0_reg\[24\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_252_1046 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_217_1166 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_197_346 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24785_ VGND VPWR VPWR VGND clk _01278_ reset_n keymem.key_mem\[6\]\[10\] sky130_fd_sc_hd__dfrtp_2
X_21997_ VPWR VGND keymem.key_mem\[3\]\[62\] _06479_ _06469_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_233_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_322 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11750_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[10\] dec_new_block\[42\]
+ _07439_ sky130_fd_sc_hd__mux2_2
XFILLER_0_212_188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23736_ keymem.prev_key0_reg\[92\] clk _00233_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20948_ VPWR VGND keymem.key_mem\[7\]\[83\] _05921_ _05899_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_230_1344 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_90_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11681_ VGND VPWR result[7] _07404_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23667_ keymem.prev_key0_reg\[23\] clk _00164_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20879_ VPWR VGND keymem.key_mem\[7\]\[51\] _05884_ _05856_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_14_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25406_ VGND VPWR VPWR VGND clk _01899_ reset_n keymem.key_mem\[2\]\[119\] sky130_fd_sc_hd__dfrtp_2
X_13420_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[125\] _07722_ keymem.key_mem\[8\]\[125\]
+ _07541_ _08898_ sky130_fd_sc_hd__a22o_2
XFILLER_0_64_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22618_ VPWR VGND VGND VPWR _06778_ keymem.key_mem_we _02708_ sky130_fd_sc_hd__nand2_2
XFILLER_0_165_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23598_ VGND VPWR VPWR VGND clk _00099_ reset_n keymem.key_mem\[14\]\[87\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_88_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25337_ VGND VPWR VPWR VGND clk _01830_ reset_n keymem.key_mem\[2\]\[50\] sky130_fd_sc_hd__dfrtp_2
X_13351_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[118\] _07702_ keymem.key_mem\[14\]\[118\]
+ _07744_ _08836_ sky130_fd_sc_hd__a22o_2
XFILLER_0_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22549_ VGND VPWR _06761_ _03287_ _01983_ _06756_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_88_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12302_ VGND VPWR VGND VPWR _07734_ keymem.key_mem\[4\]\[18\] _07884_ _07886_ _07887_
+ _07616_ sky130_fd_sc_hd__a2111o_2
X_16070_ VPWR VGND VGND VPWR _11482_ _11380_ _11375_ _11246_ _11525_ _11524_ sky130_fd_sc_hd__o221a_2
XFILLER_0_263_1164 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13282_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[111\] _07583_ keymem.key_mem\[6\]\[111\]
+ _07565_ _08774_ sky130_fd_sc_hd__a22o_2
X_25268_ VGND VPWR VPWR VGND clk _01761_ reset_n keymem.key_mem\[3\]\[109\] sky130_fd_sc_hd__dfrtp_2
X_15021_ VGND VPWR _10485_ _10446_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_60_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24219_ VGND VPWR VPWR VGND clk _00712_ reset_n keymem.key_mem\[11\]\[84\] sky130_fd_sc_hd__dfrtp_2
X_12233_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[13\] _07564_ keymem.key_mem\[2\]\[13\]
+ _07545_ _07823_ sky130_fd_sc_hd__a22o_2
X_25199_ VGND VPWR VPWR VGND clk _01692_ reset_n keymem.key_mem\[3\]\[40\] sky130_fd_sc_hd__dfrtp_2
X_12164_ VGND VPWR _07759_ _07564_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_208_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12095_ VGND VPWR _07693_ _07692_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16972_ VGND VPWR _00067_ _03100_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19760_ VGND VPWR _00667_ _05288_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_120_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15923_ VGND VPWR _11379_ _11352_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18711_ VPWR VGND VGND VPWR _04570_ _04355_ _04569_ sky130_fd_sc_hd__nand2_2
XFILLER_0_95_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19691_ VGND VPWR _00634_ _05252_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_99_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18642_ VPWR VGND VPWR VGND _04508_ _04505_ enc_block.block_w2_reg\[21\] _04504_
+ _04509_ sky130_fd_sc_hd__a22o_2
XFILLER_0_216_472 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15854_ VGND VPWR VGND VPWR _11308_ _11298_ _11250_ _11295_ _11310_ sky130_fd_sc_hd__a31o_2
XFILLER_0_235_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_494 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_235_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14805_ VGND VPWR VGND VPWR key[6] _09930_ _10270_ _10269_ _10271_ sky130_fd_sc_hd__o22a_2
XFILLER_0_207_60 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18573_ VPWR VGND VGND VPWR _04447_ _04443_ _04445_ sky130_fd_sc_hd__nand2_2
X_15785_ VGND VPWR _11241_ _11240_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12997_ VGND VPWR VGND VPWR _07808_ keymem.key_mem\[12\]\[83\] _08514_ _08516_ _08517_
+ _08480_ sky130_fd_sc_hd__a2111o_2
X_17524_ VPWR VGND VPWR VGND _03591_ _03494_ _03588_ key[244] _03527_ _03592_ sky130_fd_sc_hd__a221o_2
XFILLER_0_59_547 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14736_ VGND VPWR VGND VPWR _09945_ _09184_ _10202_ _09969_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_203_199 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11948_ VGND VPWR _07551_ _07550_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_709 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_1096 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17455_ VPWR VGND VPWR VGND _03532_ _03494_ _03529_ key[234] _03527_ _03533_ sky130_fd_sc_hd__a221o_2
X_14667_ VGND VPWR VGND VPWR _09747_ _10134_ _10129_ _10131_ _10133_ sky130_fd_sc_hd__nand4b_2
XFILLER_0_7_806 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11879_ VGND VPWR result[106] _07503_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16406_ VPWR VGND VGND VPWR _11386_ _11464_ _11469_ _11306_ _02568_ _02567_ sky130_fd_sc_hd__o221a_2
X_13618_ VGND VPWR _09090_ _09089_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17386_ VGND VPWR VGND VPWR _03473_ _03470_ _03469_ _09637_ _03472_ _09931_ sky130_fd_sc_hd__a32o_2
X_14598_ VPWR VGND VGND VPWR _09312_ _09476_ _10066_ _09423_ _09444_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_171_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_77_2_Right_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_237_Left_504 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19125_ VGND VPWR VGND VPWR _04918_ keymem.key_mem_we _02839_ _04908_ _00402_ sky130_fd_sc_hd__a31o_2
X_16337_ VPWR VGND VPWR VGND _02364_ _02420_ _02349_ _02499_ _02500_ sky130_fd_sc_hd__or4_2
X_13549_ VPWR VGND VGND VPWR enc_block.sword_ctr_reg\[1\] _09021_ enc_block.sword_ctr_reg\[0\]
+ sky130_fd_sc_hd__nor2_2
XFILLER_0_15_639 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_67_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19056_ VGND VPWR _04880_ _04879_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16268_ VPWR VGND VGND VPWR _11252_ _11385_ _02432_ _11204_ _11420_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_14_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_246_1373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_67_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18007_ VGND VPWR VGND VPWR _03736_ keymem.prev_key0_reg\[125\] _03936_ _00266_ sky130_fd_sc_hd__a21o_2
X_15219_ VGND VPWR VPWR VGND _10463_ _10464_ _10483_ _10682_ sky130_fd_sc_hd__or3_2
XFILLER_0_129_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_112_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16199_ VPWR VGND VGND VPWR _11376_ _11396_ _02364_ _11370_ _11311_ _11399_ sky130_fd_sc_hd__o32ai_2
XFILLER_0_112_368 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_103_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19958_ VGND VPWR VPWR VGND _05389_ _10099_ keymem.key_mem\[10\]\[4\] _05394_ sky130_fd_sc_hd__mux2_2
XFILLER_0_177_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_246_Left_513 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_208_951 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18909_ _04747_ _04749_ _04560_ _04748_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_78_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19889_ VGND VPWR VPWR VGND _05350_ keymem.key_mem\[11\]\[101\] _03499_ _05356_ sky130_fd_sc_hd__mux2_2
X_21920_ VGND VPWR VGND VPWR _06437_ keymem.key_mem_we _02743_ _06432_ _01678_ sky130_fd_sc_hd__a31o_2
XFILLER_0_78_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_39_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_965 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_222_442 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21851_ VGND VPWR VPWR VGND _06388_ _03654_ keymem.key_mem\[4\]\[125\] _06398_ sky130_fd_sc_hd__mux2_2
XFILLER_0_175_1191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_218_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_795 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_253_1388 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20802_ VGND VPWR VGND VPWR _05842_ keymem.key_mem_we _11149_ _05838_ _01155_ sky130_fd_sc_hd__a31o_2
X_24570_ VGND VPWR VPWR VGND clk _01063_ reset_n keymem.key_mem\[8\]\[51\] sky130_fd_sc_hd__dfrtp_2
X_21782_ VGND VPWR VPWR VGND _06355_ _03434_ keymem.key_mem\[4\]\[92\] _06362_ sky130_fd_sc_hd__mux2_2
XFILLER_0_37_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23521_ VGND VPWR VPWR VGND clk _00022_ reset_n keymem.key_mem\[14\]\[10\] sky130_fd_sc_hd__dfrtp_2
X_20733_ VGND VPWR VPWR VGND _05794_ _03580_ keymem.key_mem\[8\]\[114\] _05803_ sky130_fd_sc_hd__mux2_2
XFILLER_0_11_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_255_Left_522 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_149_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23452_ VPWR VGND VPWR VGND _07317_ _03950_ _07316_ enc_block.block_w3_reg\[25\]
+ _07126_ _02330_ sky130_fd_sc_hd__a221o_2
X_20664_ VGND VPWR VPWR VGND _05761_ _03339_ keymem.key_mem\[8\]\[81\] _05767_ sky130_fd_sc_hd__mux2_2
XFILLER_0_46_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_188_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_198 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1416 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22403_ VGND VPWR VPWR VGND _06553_ _03661_ keymem.key_mem\[2\]\[126\] _06693_ sky130_fd_sc_hd__mux2_2
XFILLER_0_149_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23383_ VGND VPWR _07256_ enc_block.block_w2_reg\[2\] enc_block.block_w0_reg\[17\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20595_ VGND VPWR VPWR VGND _05725_ _03035_ keymem.key_mem\[8\]\[48\] _05731_ sky130_fd_sc_hd__mux2_2
XFILLER_0_85_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25122_ VGND VPWR VPWR VGND clk _01615_ reset_n keymem.key_mem\[4\]\[91\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_162_279 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_60_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22334_ VGND VPWR VPWR VGND _06647_ _03443_ keymem.key_mem\[2\]\[93\] _06657_ sky130_fd_sc_hd__mux2_2
XFILLER_0_103_302 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_225_1446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_60_266 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_981 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_130_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22265_ VGND VPWR VPWR VGND _06611_ _03149_ keymem.key_mem\[2\]\[60\] _06621_ sky130_fd_sc_hd__mux2_2
XFILLER_0_225_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25053_ VGND VPWR VPWR VGND clk _01546_ reset_n keymem.key_mem\[4\]\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_170_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21216_ VGND VPWR _01349_ _06062_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24004_ VGND VPWR VPWR VGND clk _00497_ reset_n keymem.key_mem\[13\]\[125\] sky130_fd_sc_hd__dfrtp_2
X_22196_ VGND VPWR VPWR VGND _06578_ _02764_ keymem.key_mem\[2\]\[27\] _06585_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_264_Left_531 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_228_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21147_ VGND VPWR _01316_ _06026_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_22_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21078_ VGND VPWR _01283_ _05990_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_156_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_191_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20029_ VGND VPWR _00793_ _05431_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12920_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[75\] _08259_ _08447_ _08443_ _08448_
+ sky130_fd_sc_hd__o22a_2
X_24906_ VGND VPWR VPWR VGND clk _01399_ reset_n keymem.key_mem\[5\]\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_1003 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_123_1_Right_724 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_236_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24837_ VGND VPWR VPWR VGND clk _01330_ reset_n keymem.key_mem\[6\]\[62\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_214_976 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12851_ VGND VPWR enc_block.round_key\[68\] _08385_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_1058 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11802_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[4\] dec_new_block\[68\]
+ _07465_ sky130_fd_sc_hd__mux2_2
XFILLER_0_154_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_333 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15570_ VGND VPWR VGND VPWR key[13] _09930_ _11028_ _11027_ _11029_ sky130_fd_sc_hd__o22a_2
XFILLER_0_185_316 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12782_ VGND VPWR enc_block.round_key\[61\] _08323_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24768_ VGND VPWR VPWR VGND clk _01261_ reset_n keymem.key_mem\[7\]\[121\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_68_355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_90_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14521_ VPWR VGND VGND VPWR _09990_ _09989_ _09986_ _09931_ _09930_ key[3] sky130_fd_sc_hd__o2111a_2
X_11733_ VGND VPWR result[33] _07430_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_68_377 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23719_ keymem.prev_key0_reg\[75\] clk _00216_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_3_1001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24699_ VGND VPWR VPWR VGND clk _01192_ reset_n keymem.key_mem\[7\]\[52\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_51_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17240_ VPWR VGND VGND VPWR _08936_ _03342_ key[82] sky130_fd_sc_hd__nor2_2
X_14452_ VPWR VGND VPWR VGND _09591_ _09920_ _09592_ _09590_ _09921_ sky130_fd_sc_hd__or4_2
XFILLER_0_3_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11664_ VGND VPWR VPWR VGND encdec _07396_ next sky130_fd_sc_hd__and2b_2
XFILLER_0_193_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13403_ VGND VPWR VGND VPWR _07838_ keymem.key_mem\[11\]\[123\] _08878_ _08880_ _08883_
+ _08882_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_3_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17171_ VGND VPWR _03280_ _09541_ _00086_ _03279_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_14383_ VGND VPWR VGND VPWR _09852_ _09851_ _09853_ keymem.prev_key0_reg\[98\] sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_1121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_144_1_Left_411 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16122_ VPWR VGND VGND VPWR _11404_ _11236_ _11375_ _11298_ _11576_ _11575_ sky130_fd_sc_hd__o221a_2
X_13334_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[116\] _08714_ _08820_ _08814_ _08821_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_243_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_789 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16053_ VGND VPWR VGND VPWR _11508_ _11273_ _11289_ _11227_ _11226_ sky130_fd_sc_hd__and4_2
X_13265_ VGND VPWR VGND VPWR _08759_ _08008_ keymem.key_mem\[2\]\[109\] _08756_ _08758_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_267_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_631 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_32_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15004_ VPWR VGND VPWR VGND _10456_ _10435_ _10429_ _10419_ _10468_ sky130_fd_sc_hd__or4_2
XFILLER_0_122_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12216_ VGND VPWR _07807_ _07806_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_62_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_267_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13196_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[103\] _07782_ keymem.key_mem\[6\]\[103\]
+ _07739_ _08696_ sky130_fd_sc_hd__a22o_2
XFILLER_0_161_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19812_ VGND VPWR VPWR VGND _05314_ keymem.key_mem\[11\]\[64\] _03194_ _05316_ sky130_fd_sc_hd__mux2_2
XFILLER_0_202_1243 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12147_ VGND VPWR _07743_ _07742_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_264_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19743_ VGND VPWR _00659_ _05279_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16955_ VGND VPWR _00065_ _03085_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_263_364 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_208_269 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12078_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[3\] _07645_ _07677_ _07664_ _07678_
+ sky130_fd_sc_hd__o22a_2
X_15906_ VGND VPWR VGND VPWR _11262_ _11282_ _11361_ _11318_ _11362_ sky130_fd_sc_hd__o22a_2
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16886_ VGND VPWR VPWR VGND _03020_ _11110_ _03023_ _03022_ _03021_ sky130_fd_sc_hd__o211a_2
X_19674_ VPWR VGND VGND VPWR _05242_ _05240_ _05241_ sky130_fd_sc_hd__nand2_2
XFILLER_0_154_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15837_ VGND VPWR VGND VPWR _11293_ _11291_ _11290_ _11224_ _11292_ _11287_ sky130_fd_sc_hd__a32o_2
X_18625_ VPWR VGND _04494_ _04493_ enc_block.round_key\[83\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_188_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_188_154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_151_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15768_ VGND VPWR _11224_ _11223_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18556_ VPWR VGND _04432_ _04431_ enc_block.round_key\[76\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_249_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_133_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14719_ VGND VPWR VPWR VGND keymem.round_ctr_reg\[0\] _10185_ _10141_ _10186_ sky130_fd_sc_hd__mux2_2
X_17507_ VPWR VGND VGND VPWR _03577_ key[242] _09868_ sky130_fd_sc_hd__nand2_2
XFILLER_0_59_388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18487_ VPWR VGND _04370_ _04369_ enc_block.round_key\[69\] VPWR VGND sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_107_2_Left_578 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_170_13 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15699_ VGND VPWR VPWR VGND _11155_ keymem.prev_key1_reg\[80\] _11152_ _11153_ _09729_
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_30_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_200_670 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_191_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17438_ VPWR VGND VPWR VGND _03517_ _03494_ _03513_ key[232] _03366_ _03518_ sky130_fd_sc_hd__a221o_2
XFILLER_0_16_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_1_Left_343 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_144_224 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_55_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17369_ VGND VPWR VPWR VGND _10323_ key[223] _03458_ _10281_ _03457_ sky130_fd_sc_hd__o211a_2
X_19108_ VGND VPWR VGND VPWR _04909_ keymem.key_mem_we _02608_ _04908_ _00394_ sky130_fd_sc_hd__a31o_2
XFILLER_0_28_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20380_ VGND VPWR _05617_ _03279_ _00958_ _05532_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_179_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_183_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19039_ VGND VPWR VGND VPWR _03959_ block[62] _04865_ _04864_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_24_981 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_169_2_Left_640 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_288 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22050_ VPWR VGND keymem.key_mem\[3\]\[87\] _06507_ _06484_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_80_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_140_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_144_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21001_ VGND VPWR _01248_ _05948_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_56_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_697 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_142_1190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_887 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_195_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_39_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25740_ keymem.prev_key1_reg\[56\] clk _02233_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22952_ VGND VPWR VGND VPWR _02209_ _06938_ _06916_ keymem.prev_key1_reg\[32\] sky130_fd_sc_hd__o21a_2
XFILLER_0_128_92 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_39_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21903_ VGND VPWR VGND VPWR _06428_ keymem.key_mem_we _02340_ _06420_ _01670_ sky130_fd_sc_hd__a31o_2
XFILLER_0_190_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25671_ VGND VPWR VPWR VGND clk _02164_ reset_n keymem.rcon_reg\[0\] sky130_fd_sc_hd__dfrtp_2
X_22883_ VGND VPWR VPWR VGND _06878_ _06895_ keymem.prev_key1_reg\[6\] _06896_ sky130_fd_sc_hd__mux2_2
XFILLER_0_214_1114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_151_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24622_ VGND VPWR VPWR VGND clk _01115_ reset_n keymem.key_mem\[8\]\[103\] sky130_fd_sc_hd__dfrtp_2
X_21834_ VGND VPWR _01640_ _06389_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_190_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_194_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_151_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_467 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24553_ VGND VPWR VPWR VGND clk _01046_ reset_n keymem.key_mem\[8\]\[34\] sky130_fd_sc_hd__dfrtp_2
X_21765_ VGND VPWR VPWR VGND _06344_ _03364_ keymem.key_mem\[4\]\[84\] _06353_ sky130_fd_sc_hd__mux2_2
X_23504_ VGND VPWR _04301_ _07362_ _07364_ _07363_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_20716_ VGND VPWR _05794_ _05675_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_4_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24484_ VGND VPWR VPWR VGND clk _00977_ reset_n keymem.key_mem\[9\]\[93\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_135_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21696_ VGND VPWR VPWR VGND _06308_ _03067_ keymem.key_mem\[4\]\[51\] _06317_ sky130_fd_sc_hd__mux2_2
XFILLER_0_149_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_110_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_190_330 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23435_ VPWR VGND VPWR VGND _07302_ block[23] _04139_ enc_block.block_w0_reg\[23\]
+ _04138_ _07303_ sky130_fd_sc_hd__a221o_2
XFILLER_0_19_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20647_ VGND VPWR VPWR VGND _05747_ _03267_ keymem.key_mem\[8\]\[73\] _05758_ sky130_fd_sc_hd__mux2_2
XFILLER_0_184_1268 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23366_ VPWR VGND VGND VPWR _07241_ enc_block.block_w0_reg\[23\] _07239_ sky130_fd_sc_hd__nand2_2
X_20578_ VGND VPWR VPWR VGND _05714_ _02955_ keymem.key_mem\[8\]\[40\] _05722_ sky130_fd_sc_hd__mux2_2
XFILLER_0_184_1279 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_150_238 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25105_ VGND VPWR VPWR VGND clk _01598_ reset_n keymem.key_mem\[4\]\[74\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_150_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22317_ VGND VPWR _01864_ _06648_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_428 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_225_1254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23297_ VPWR VGND VGND VPWR _07179_ _07175_ _07177_ sky130_fd_sc_hd__nand2_2
XFILLER_0_103_143 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_162_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_951 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13050_ VPWR VGND VPWR VGND _08564_ keymem.key_mem\[10\]\[88\] _07876_ keymem.key_mem\[12\]\[88\]
+ _07894_ _08565_ sky130_fd_sc_hd__a221o_2
X_25036_ VGND VPWR VPWR VGND clk _01529_ reset_n keymem.key_mem\[4\]\[5\] sky130_fd_sc_hd__dfrtp_2
X_22248_ VGND VPWR _01831_ _06612_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_44_1062 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12001_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[0\] _07603_ keymem.key_mem\[11\]\[0\]
+ _07600_ _07604_ sky130_fd_sc_hd__a22o_2
X_22179_ VGND VPWR VPWR VGND _06565_ _02409_ keymem.key_mem\[2\]\[19\] _06576_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_90_2_Left_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_108_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16740_ VGND VPWR VGND VPWR _02890_ _09721_ _09795_ key[34] sky130_fd_sc_hd__o21a_2
X_13952_ VGND VPWR VGND VPWR _09350_ _09419_ _09423_ _09420_ _09424_ sky130_fd_sc_hd__o22a_2
XFILLER_0_57_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_868 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12903_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[74\] _07649_ keymem.key_mem\[9\]\[74\]
+ _07716_ _08432_ sky130_fd_sc_hd__a22o_2
X_16671_ VGND VPWR _02825_ keymem.prev_key0_reg\[30\] _02824_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_13883_ VGND VPWR _09355_ _09354_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_202_913 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_124_1_Right_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15622_ VPWR VGND VPWR VGND _11080_ _10865_ _11079_ sky130_fd_sc_hd__or2_2
X_18410_ VPWR VGND VPWR VGND _04301_ _08940_ _10316_ sky130_fd_sc_hd__or2_2
X_12834_ VPWR VGND VPWR VGND _08369_ keymem.key_mem\[5\]\[67\] _07613_ keymem.key_mem\[8\]\[67\]
+ _07903_ _08370_ sky130_fd_sc_hd__a221o_2
X_19390_ VGND VPWR VPWR VGND _04876_ _05087_ keymem.key_mem\[13\]\[126\] _05088_ sky130_fd_sc_hd__mux2_2
XFILLER_0_33_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18341_ VPWR VGND _04239_ _04238_ enc_block.round_key\[120\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15553_ VPWR VGND VPWR VGND _10694_ _10807_ _11011_ _10624_ _11012_ sky130_fd_sc_hd__or4_2
XFILLER_0_51_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12765_ VPWR VGND VPWR VGND _08307_ keymem.key_mem\[8\]\[60\] _08211_ keymem.key_mem\[1\]\[60\]
+ _07715_ _08308_ sky130_fd_sc_hd__a221o_2
X_14504_ VGND VPWR VGND VPWR _09693_ _09047_ _09087_ _09061_ _09973_ sky130_fd_sc_hd__a31o_2
XFILLER_0_173_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11716_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[25\] dec_new_block\[25\]
+ _07422_ sky130_fd_sc_hd__mux2_2
X_18272_ _04174_ _04176_ _04008_ _04175_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_166_360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15484_ VGND VPWR VPWR VGND _10457_ _10430_ _10443_ _10944_ sky130_fd_sc_hd__or3_2
XFILLER_0_83_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12696_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[53\] _07583_ keymem.key_mem\[11\]\[53\]
+ _07861_ _08246_ sky130_fd_sc_hd__a22o_2
X_17223_ VPWR VGND VPWR VGND _03327_ keymem.prev_key0_reg\[80\] _09517_ _11441_ _03326_
+ _09513_ sky130_fd_sc_hd__o311a_2
X_14435_ VPWR VGND VPWR VGND _09568_ _09593_ _09569_ _09903_ _09904_ sky130_fd_sc_hd__or4_2
XFILLER_0_181_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_126_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11647_ VPWR VGND VPWR VGND _07384_ keymem.ready_new sky130_fd_sc_hd__inv_2
XFILLER_0_4_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17154_ VPWR VGND VPWR VGND _03265_ _03263_ _09517_ _02957_ _03264_ _09513_ sky130_fd_sc_hd__o311a_2
X_14366_ VPWR VGND VGND VPWR _09103_ _09146_ _09127_ _09211_ _09836_ _09835_ sky130_fd_sc_hd__o221a_2
XFILLER_0_68_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16105_ VGND VPWR VPWR VGND _11558_ _11552_ _11549_ _11559_ sky130_fd_sc_hd__mux2_2
X_13317_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[115\] _07812_ keymem.key_mem\[9\]\[115\]
+ _07716_ _08805_ sky130_fd_sc_hd__a22o_2
X_17085_ VGND VPWR _00077_ _03203_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14297_ VGND VPWR VGND VPWR _09323_ _09332_ _09366_ _09363_ _09754_ _09767_ sky130_fd_sc_hd__o32a_2
XFILLER_0_29_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16036_ VPWR VGND VGND VPWR _11280_ _11491_ _11284_ sky130_fd_sc_hd__nor2_2
X_13248_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[108\] _07652_ keymem.key_mem\[9\]\[108\]
+ _07717_ _08743_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_237_832 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13179_ VGND VPWR VGND VPWR _07908_ keymem.key_mem\[6\]\[101\] _08678_ _08680_ _08681_
+ _08599_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_199_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17987_ VGND VPWR VPWR VGND _03281_ key[247] keymem.prev_key1_reg\[119\] _03923_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_209_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_165_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19726_ VGND VPWR VPWR VGND _05270_ keymem.key_mem\[11\]\[23\] _02661_ _05271_ sky130_fd_sc_hd__mux2_2
XFILLER_0_139_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16938_ VGND VPWR VGND VPWR _02464_ _02342_ _03070_ _02463_ sky130_fd_sc_hd__nand3_2
XPHY_EDGE_ROW_239_Right_108 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_215_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19657_ VGND VPWR _00620_ _05232_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_40_Left_308 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16869_ VGND VPWR _00057_ _03007_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_219_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_220_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18608_ VGND VPWR _04478_ _03965_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19588_ VGND VPWR VGND VPWR _05196_ keymem.key_mem_we _03393_ _05187_ _00587_ sky130_fd_sc_hd__a31o_2
XFILLER_0_172_1183 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_133_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18539_ VGND VPWR _04416_ enc_block.block_w3_reg\[10\] enc_block.block_w3_reg\[15\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21550_ VGND VPWR VPWR VGND _06231_ _03560_ keymem.key_mem\[5\]\[111\] _06239_ sky130_fd_sc_hd__mux2_2
XFILLER_0_34_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_138 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_23_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_7_444 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_56_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20501_ VGND VPWR VPWR VGND _05680_ _09991_ keymem.key_mem\[8\]\[3\] _05682_ sky130_fd_sc_hd__mux2_2
XFILLER_0_117_246 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21481_ VGND VPWR VPWR VGND _06196_ _03314_ keymem.key_mem\[5\]\[78\] _06203_ sky130_fd_sc_hd__mux2_2
XFILLER_0_1_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_257 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_745 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_99_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23220_ VGND VPWR _07109_ enc_block.block_w3_reg\[25\] enc_block.block_w3_reg\[26\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20432_ VGND VPWR _00983_ _05644_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_132_216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_226_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23151_ VGND VPWR VPWR VGND _07054_ _07059_ keymem.prev_key1_reg\[110\] _07060_ sky130_fd_sc_hd__mux2_2
X_20363_ VGND VPWR _00950_ _05608_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_259_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22102_ VGND VPWR VPWR VGND _06527_ _05058_ keymem.key_mem\[3\]\[112\] _06534_ sky130_fd_sc_hd__mux2_2
X_23082_ VGND VPWR VGND VPWR _02261_ _07016_ _07010_ keymem.prev_key1_reg\[84\] sky130_fd_sc_hd__o21a_2
XFILLER_0_144_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20294_ VGND VPWR _00917_ _05572_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_247_629 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_80_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22033_ VGND VPWR _06498_ _06403_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_45_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_197_Left_464 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_80 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_254_172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_199_216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23984_ VGND VPWR VPWR VGND clk _00477_ reset_n keymem.key_mem\[13\]\[105\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_242_356 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_39_1131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25723_ keymem.prev_key1_reg\[39\] clk _02216_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_225_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22935_ VGND VPWR _06928_ _10085_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_97_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25654_ VGND VPWR VPWR VGND clk _02147_ reset_n keymem.key_mem\[0\]\[111\] sky130_fd_sc_hd__dfrtp_2
X_22866_ VGND VPWR _06884_ _06883_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_151_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1283 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24605_ VGND VPWR VPWR VGND clk _01098_ reset_n keymem.key_mem\[8\]\[86\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_112_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21817_ VGND VPWR _01632_ _06380_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_91_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25585_ VGND VPWR VPWR VGND clk _02078_ reset_n keymem.key_mem\[0\]\[42\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_151_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22797_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[100\] _06850_ _06849_ _05033_ _02136_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_241_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12550_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[39\] _07893_ _08113_ _08109_ _08114_
+ sky130_fd_sc_hd__o22a_2
X_24536_ VGND VPWR VPWR VGND clk _01029_ reset_n keymem.key_mem\[8\]\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21748_ VGND VPWR _06344_ _06262_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_52_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_4_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_328 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_65_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24467_ VGND VPWR VPWR VGND clk _00960_ reset_n keymem.key_mem\[9\]\[76\] sky130_fd_sc_hd__dfrtp_2
X_12481_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[33\] _07924_ keymem.key_mem\[2\]\[33\]
+ _07816_ _08051_ sky130_fd_sc_hd__a22o_2
X_21679_ VGND VPWR _06308_ _06262_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14220_ VGND VPWR VGND VPWR _09113_ _09109_ _09125_ _09160_ _09691_ sky130_fd_sc_hd__o22a_2
X_23418_ VPWR VGND VPWR VGND _07287_ block[21] _04139_ enc_block.block_w0_reg\[21\]
+ _04138_ _07288_ sky130_fd_sc_hd__a221o_2
XFILLER_0_190_171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24398_ VGND VPWR VPWR VGND clk _00891_ reset_n keymem.key_mem\[9\]\[7\] sky130_fd_sc_hd__dfrtp_2
X_14151_ VPWR VGND VPWR VGND _09261_ _09245_ _09314_ _09254_ _09622_ sky130_fd_sc_hd__or4_2
XFILLER_0_22_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23349_ _07224_ _07226_ _03982_ _07225_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_85_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13102_ VPWR VGND VPWR VGND _08611_ keymem.key_mem\[3\]\[93\] _08009_ keymem.key_mem\[8\]\[93\]
+ _08265_ _08612_ sky130_fd_sc_hd__a221o_2
XFILLER_0_46_1168 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_162_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14082_ VGND VPWR VGND VPWR _09553_ _09291_ _09339_ _09307_ _09306_ sky130_fd_sc_hd__and4_2
XFILLER_0_131_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_123_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13033_ VGND VPWR enc_block.round_key\[86\] _08549_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25019_ VGND VPWR VPWR VGND clk _01512_ reset_n keymem.key_mem\[5\]\[116\] sky130_fd_sc_hd__dfrtp_2
X_17910_ VGND VPWR VGND VPWR _03730_ keymem.prev_key0_reg\[94\] _03870_ _03450_ _00235_
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_63_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18890_ VGND VPWR VGND VPWR _04732_ _04505_ _04731_ _04730_ sky130_fd_sc_hd__o21a_2
XFILLER_0_28_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17841_ VGND VPWR VPWR VGND _03814_ _03823_ keymem.prev_key0_reg\[72\] _03824_ sky130_fd_sc_hd__mux2_2
X_14984_ VPWR VGND VPWR VGND _10447_ _10409_ _10403_ _10439_ _10448_ sky130_fd_sc_hd__or4_2
X_17772_ VGND VPWR _03777_ _03674_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19511_ VGND VPWR VGND VPWR _05155_ keymem.key_mem_we _03068_ _05135_ _00551_ sky130_fd_sc_hd__a31o_2
XPHY_EDGE_ROW_201_Left_468 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_156_1145 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13935_ VGND VPWR VPWR VGND _09304_ _09315_ _09297_ _09407_ sky130_fd_sc_hd__or3_2
X_16723_ VGND VPWR _00044_ _02874_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19442_ VGND VPWR VGND VPWR _05118_ keymem.key_mem_we _02410_ _05109_ _00519_ sky130_fd_sc_hd__a31o_2
X_16654_ VPWR VGND VGND VPWR _02808_ _02809_ keylen sky130_fd_sc_hd__nor2_2
X_13866_ VGND VPWR _09338_ _09337_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_125_1_Right_726 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_134_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15605_ VGND VPWR VGND VPWR _10458_ _10592_ _10524_ _10611_ _11063_ sky130_fd_sc_hd__o22a_2
XFILLER_0_201_242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12817_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[65\] _07578_ keymem.key_mem\[1\]\[65\]
+ _07855_ _08355_ sky130_fd_sc_hd__a22o_2
XFILLER_0_9_709 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_130_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19373_ VGND VPWR _00492_ _05076_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16585_ VGND VPWR _02743_ _02742_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13797_ VGND VPWR _09269_ _08944_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_134_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_151_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15536_ VPWR VGND VPWR VGND _10650_ _10621_ _10941_ _10994_ _10995_ sky130_fd_sc_hd__or4bb_2
X_18324_ VPWR VGND VGND VPWR _04223_ _04224_ _04190_ sky130_fd_sc_hd__nor2_2
XFILLER_0_70_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12748_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[58\] _07759_ keymem.key_mem\[12\]\[58\]
+ _07673_ _08293_ sky130_fd_sc_hd__a22o_2
XFILLER_0_139_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_44_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18255_ VPWR VGND VPWR VGND _04160_ _04040_ _04158_ enc_block.block_w0_reg\[16\]
+ _04097_ _00290_ sky130_fd_sc_hd__a221o_2
X_15467_ VPWR VGND VGND VPWR _10639_ _10927_ _10593_ sky130_fd_sc_hd__nor2_2
XFILLER_0_71_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12679_ VGND VPWR enc_block.round_key\[51\] _08230_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17206_ VGND VPWR VPWR VGND _03311_ _03312_ keymem.prev_key0_reg\[78\] _10327_ _11092_
+ sky130_fd_sc_hd__a31oi_2
XPHY_EDGE_ROW_210_Left_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14418_ VGND VPWR VGND VPWR _09448_ _09447_ _09885_ _09473_ _09887_ _09886_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_4_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_114_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18186_ VGND VPWR _04097_ _03974_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15398_ VGND VPWR VGND VPWR _10701_ _10858_ _10859_ _10699_ _10702_ sky130_fd_sc_hd__nor4_2
XFILLER_0_245_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17137_ VGND VPWR VPWR VGND _02936_ keymem.prev_key0_reg\[71\] _03250_ _03249_ _03248_
+ sky130_fd_sc_hd__o211a_2
X_14349_ VGND VPWR VGND VPWR _09122_ _09100_ _09687_ _09141_ _09819_ sky130_fd_sc_hd__o22a_2
XFILLER_0_64_1257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_141_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17068_ VGND VPWR VPWR VGND _03187_ _09530_ _03188_ _09529_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_180_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_578 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_21_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16019_ VPWR VGND VPWR VGND _11473_ _11306_ _11325_ _11286_ _11338_ _11474_ sky130_fd_sc_hd__a221o_2
XFILLER_0_141_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_85_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_23 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_85_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_243_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_221_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_250_Right_119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_178_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1028 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_109_83 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19709_ VGND VPWR VPWR VGND _05259_ keymem.key_mem\[11\]\[15\] _11149_ _05262_ sky130_fd_sc_hd__mux2_2
XFILLER_0_197_709 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_174_1245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_251_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20981_ VGND VPWR VPWR VGND _05934_ _05031_ keymem.key_mem\[7\]\[99\] _05938_ sky130_fd_sc_hd__mux2_2
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22720_ VGND VPWR _02090_ _06825_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_251_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_149_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_152_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_82 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22651_ VGND VPWR _02050_ _06796_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_113_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21602_ VGND VPWR VPWR VGND _06263_ _10283_ keymem.key_mem\[4\]\[6\] _06268_ sky130_fd_sc_hd__mux2_2
X_25370_ VGND VPWR VPWR VGND clk _01863_ reset_n keymem.key_mem\[2\]\[83\] sky130_fd_sc_hd__dfrtp_2
X_22582_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[96\] _06767_ _06766_ _05024_ _02004_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_164_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24321_ VGND VPWR VPWR VGND clk _00814_ reset_n keymem.key_mem\[10\]\[58\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21533_ VGND VPWR VPWR VGND _06220_ _03511_ keymem.key_mem\[5\]\[103\] _06230_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_520 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_141_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24252_ VGND VPWR VPWR VGND clk _00745_ reset_n keymem.key_mem\[11\]\[117\] sky130_fd_sc_hd__dfrtp_2
X_21464_ VGND VPWR VPWR VGND _06184_ _03245_ keymem.key_mem\[5\]\[70\] _06194_ sky130_fd_sc_hd__mux2_2
XFILLER_0_263_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_160_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23203_ VGND VPWR VPWR VGND _07093_ enc_block.block_w3_reg\[0\] _03971_ _07094_ sky130_fd_sc_hd__mux2_2
X_20415_ VGND VPWR _00975_ _05635_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24183_ VGND VPWR VPWR VGND clk _00676_ reset_n keymem.key_mem\[11\]\[48\] sky130_fd_sc_hd__dfrtp_2
X_21395_ VGND VPWR VPWR VGND _06151_ _02923_ keymem.key_mem\[5\]\[37\] _06158_ sky130_fd_sc_hd__mux2_2
XFILLER_0_181_1249 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_4_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23134_ VGND VPWR VGND VPWR _03521_ _03520_ _03524_ _07048_ sky130_fd_sc_hd__a21o_2
X_20346_ VGND VPWR _00942_ _05599_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_113_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23065_ VPWR VGND VPWR VGND _03312_ _03310_ _03794_ _03309_ _07006_ sky130_fd_sc_hd__a22o_2
X_20277_ VGND VPWR _00909_ _05563_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_228_640 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22016_ VPWR VGND keymem.key_mem\[3\]\[71\] _06489_ _06484_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_200_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_179_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_216_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_168_2_Right_240 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_236_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_632 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_200_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_196_1481 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23967_ VGND VPWR VPWR VGND clk _00460_ reset_n keymem.key_mem\[13\]\[88\] sky130_fd_sc_hd__dfrtp_2
X_11981_ VGND VPWR _07584_ _07583_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_19_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_153_1_Left_420 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13720_ VGND VPWR VGND VPWR _09191_ _09059_ _09060_ _09188_ _09192_ sky130_fd_sc_hd__a31o_2
X_25706_ keymem.prev_key1_reg\[22\] clk _02199_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_242_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22918_ VGND VPWR VGND VPWR _06917_ _02468_ _06891_ _02478_ _06892_ sky130_fd_sc_hd__a211o_2
X_23898_ VGND VPWR VPWR VGND clk _00391_ reset_n keymem.key_mem\[13\]\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13651_ VPWR VGND VPWR VGND _09014_ _09005_ _08991_ _08977_ _09123_ sky130_fd_sc_hd__or4_2
X_25637_ VGND VPWR VPWR VGND clk _02130_ reset_n keymem.key_mem\[0\]\[94\] sky130_fd_sc_hd__dfrtp_2
X_22849_ VGND VPWR _02172_ _06872_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_78_280 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_239 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12602_ VGND VPWR VGND VPWR _08161_ _07703_ keymem.key_mem\[7\]\[44\] _08160_ _07746_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_196_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16370_ _11224_ _02533_ _11412_ _11292_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_17_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13582_ VGND VPWR VGND VPWR _09050_ _08999_ _09054_ _09053_ sky130_fd_sc_hd__a21oi_2
X_25568_ VGND VPWR VPWR VGND clk _02061_ reset_n keymem.key_mem\[0\]\[25\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15321_ VGND VPWR VGND VPWR _10485_ _10519_ _10498_ _10546_ _10783_ sky130_fd_sc_hd__o22a_2
XFILLER_0_93_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12533_ VPWR VGND VPWR VGND _08097_ keymem.key_mem\[5\]\[38\] _08096_ keymem.key_mem\[14\]\[38\]
+ _07721_ _08098_ sky130_fd_sc_hd__a221o_2
X_24519_ VGND VPWR VPWR VGND clk _01012_ reset_n keymem.key_mem\[8\]\[0\] sky130_fd_sc_hd__dfrtp_2
X_25499_ VGND VPWR VPWR VGND clk _01992_ reset_n keymem.key_mem\[1\]\[84\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18040_ VPWR VGND _03962_ _03961_ _03960_ VPWR VGND sky130_fd_sc_hd__xor2_2
X_15252_ VGND VPWR VGND VPWR _10715_ _10572_ _10543_ _10633_ _10627_ _10714_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_136_385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_862 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12464_ VGND VPWR VGND VPWR _08036_ _07841_ keymem.key_mem\[4\]\[31\] _08033_ _08035_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_168_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_53_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_87_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_40 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_670 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14203_ VGND VPWR VGND VPWR _09674_ _09671_ _09215_ _09672_ _09673_ sky130_fd_sc_hd__a211o_2
XFILLER_0_262_1037 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15183_ VGND VPWR VGND VPWR _10572_ _10608_ _10536_ _10646_ _10580_ _10647_ sky130_fd_sc_hd__o32a_2
X_12395_ VGND VPWR VGND VPWR _07973_ _07968_ keymem.key_mem\[9\]\[25\] _07970_ _07972_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_151_366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_854 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_205_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14134_ VGND VPWR VGND VPWR _09605_ _09602_ _09248_ _09603_ _09604_ sky130_fd_sc_hd__a211o_2
XFILLER_0_22_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19991_ VGND VPWR _00775_ _05411_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_22_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18942_ VPWR VGND VGND VPWR _04778_ _04779_ _04191_ sky130_fd_sc_hd__nor2_2
XFILLER_0_201_1319 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14065_ VGND VPWR _09537_ _09536_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_24_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13016_ VPWR VGND VPWR VGND _08533_ keymem.key_mem\[13\]\[85\] _07834_ keymem.key_mem\[4\]\[85\]
+ _07914_ _08534_ sky130_fd_sc_hd__a221o_2
XFILLER_0_20_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_116_2_Left_587 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18873_ VPWR VGND VGND VPWR _04654_ _04717_ _04116_ sky130_fd_sc_hd__nor2_2
XFILLER_0_98_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_123_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17824_ VGND VPWR _00208_ _03811_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_59_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_85_1_Left_352 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_261_440 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_55_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14967_ enc_block.sword_ctr_reg\[1\] _10431_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[15\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_238_1286 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17755_ VGND VPWR _00183_ _03767_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_57_1061 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_221_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16706_ VPWR VGND VPWR VGND _02859_ key[159] _10286_ sky130_fd_sc_hd__or2_2
X_13918_ VPWR VGND VPWR VGND _09328_ _09309_ _09339_ _09306_ _09390_ sky130_fd_sc_hd__or4_2
X_17686_ VGND VPWR VPWR VGND _03703_ _03720_ keymem.prev_key0_reg\[20\] _03721_ sky130_fd_sc_hd__mux2_2
X_14898_ VGND VPWR VGND VPWR _10362_ _10361_ _10363_ keymem.prev_key0_reg\[103\] sky130_fd_sc_hd__a21oi_2
XFILLER_0_76_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_134_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19425_ VGND VPWR _05109_ _05092_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13849_ VGND VPWR VGND VPWR _09321_ _09284_ _09283_ keymem.prev_key1_reg\[29\] _08969_
+ _08964_ sky130_fd_sc_hd__a32o_2
X_16637_ VGND VPWR VGND VPWR _02791_ _10360_ _02789_ _02790_ _02792_ sky130_fd_sc_hd__a31o_2
XPHY_EDGE_ROW_126_1_Right_727 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_134_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19356_ VGND VPWR VPWR VGND _05046_ _05064_ keymem.key_mem\[13\]\[115\] _05065_ sky130_fd_sc_hd__mux2_2
X_16568_ _09759_ _02726_ keymem.round_ctr_reg\[0\] _09789_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_70_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18307_ VGND VPWR VGND VPWR _04208_ _03982_ _04207_ _04206_ sky130_fd_sc_hd__o21a_2
XFILLER_0_169_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15519_ VGND VPWR _00024_ _10978_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16499_ VPWR VGND VPWR VGND _02659_ _02649_ _02648_ key[151] _11043_ _02660_ sky130_fd_sc_hd__a221o_2
X_19287_ VPWR VGND keymem.key_mem\[13\]\[92\] _05019_ _04879_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_127_363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_723 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18238_ _04143_ _04145_ _03981_ _04144_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_66_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_142_322 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_154_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_810 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_245_1257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18169_ VPWR VGND VGND VPWR _04081_ _04082_ _04077_ sky130_fd_sc_hd__nor2_2
XFILLER_0_64_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20200_ VGND VPWR VPWR VGND _05515_ _03613_ keymem.key_mem\[10\]\[119\] _05521_ sky130_fd_sc_hd__mux2_2
XFILLER_0_25_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21180_ VGND VPWR VPWR VGND _06040_ _03193_ keymem.key_mem\[6\]\[64\] _06044_ sky130_fd_sc_hd__mux2_2
XFILLER_0_64_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_106_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_141_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20131_ VGND VPWR VPWR VGND _05482_ _03383_ keymem.key_mem\[10\]\[86\] _05485_ sky130_fd_sc_hd__mux2_2
XFILLER_0_187_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_96_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20062_ VGND VPWR VPWR VGND _05446_ _03083_ keymem.key_mem\[10\]\[53\] _05449_ sky130_fd_sc_hd__mux2_2
XFILLER_0_42_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1028 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_253_941 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24870_ VGND VPWR VPWR VGND clk _01363_ reset_n keymem.key_mem\[6\]\[95\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_224_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23821_ VGND VPWR VPWR VGND clk _00314_ reset_n enc_block.block_w1_reg\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23752_ keymem.prev_key0_reg\[108\] clk _00249_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_136_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20964_ VPWR VGND keymem.key_mem\[7\]\[91\] _05929_ _05823_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_67_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22703_ VGND VPWR _06820_ _06779_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_117_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_152_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23683_ keymem.prev_key0_reg\[39\] clk _00180_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20895_ VGND VPWR VGND VPWR _05892_ keymem.key_mem_we _03130_ _05864_ _01198_ sky130_fd_sc_hd__a31o_2
XFILLER_0_36_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25422_ VGND VPWR VPWR VGND clk _01915_ reset_n keymem.key_mem\[1\]\[7\] sky130_fd_sc_hd__dfrtp_2
X_22634_ VGND VPWR VPWR VGND _06785_ keymem.key_mem\[0\]\[6\] _10284_ _06788_ sky130_fd_sc_hd__mux2_2
XFILLER_0_152_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_113_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_1110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_64_946 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25353_ VGND VPWR VPWR VGND clk _01846_ reset_n keymem.key_mem\[2\]\[66\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_187_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22565_ VGND VPWR _06767_ _06696_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_192_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24304_ VGND VPWR VPWR VGND clk _00797_ reset_n keymem.key_mem\[10\]\[41\] sky130_fd_sc_hd__dfrtp_2
X_21516_ VGND VPWR _01490_ _06221_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_90_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25284_ VGND VPWR VPWR VGND clk _01777_ reset_n keymem.key_mem\[3\]\[125\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_873 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_84_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22496_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[46\] _06737_ _06736_ _04947_ _01954_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_263_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24235_ VGND VPWR VPWR VGND clk _00728_ reset_n keymem.key_mem\[11\]\[100\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_228_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21447_ VGND VPWR _01457_ _06185_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_160_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_43_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24166_ VGND VPWR VPWR VGND clk _00659_ reset_n keymem.key_mem\[11\]\[31\] sky130_fd_sc_hd__dfrtp_2
X_12180_ VGND VPWR VGND VPWR _07774_ _07579_ keymem.key_mem\[12\]\[9\] _07770_ _07773_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_32_887 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21378_ VGND VPWR VPWR VGND _06140_ _02811_ keymem.key_mem\[5\]\[29\] _06149_ sky130_fd_sc_hd__mux2_2
XFILLER_0_124_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23117_ VGND VPWR _02275_ _07037_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_248_746 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20329_ VGND VPWR _00934_ _05590_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24097_ VGND VPWR VPWR VGND clk _00590_ reset_n keymem.key_mem\[12\]\[90\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_198_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23048_ VPWR VGND VGND VPWR _06995_ _06996_ keylen sky130_fd_sc_hd__nor2_2
XFILLER_0_21_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_159_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_194_1418 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15870_ VPWR VGND VPWR VGND _11206_ _11229_ _11207_ _11225_ _11326_ sky130_fd_sc_hd__or4_2
XFILLER_0_95_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_654 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_169_2_Right_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_216_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14821_ VGND VPWR _10286_ _09729_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_95_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24999_ VGND VPWR VPWR VGND clk _01492_ reset_n keymem.key_mem\[5\]\[96\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_235_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14752_ VGND VPWR VGND VPWR _09113_ _09156_ _09646_ _09177_ _09040_ _10218_ sky130_fd_sc_hd__o32a_2
X_17540_ VGND VPWR VGND VPWR _03606_ _03603_ _03602_ _09637_ _03605_ _09931_ sky130_fd_sc_hd__a32o_2
XFILLER_0_263_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11964_ VGND VPWR _07567_ _07566_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13703_ VGND VPWR VGND VPWR _09174_ _09109_ _09167_ _09100_ _09175_ sky130_fd_sc_hd__o22a_2
X_17471_ VGND VPWR VPWR VGND _03029_ _03545_ key[109] _03546_ sky130_fd_sc_hd__mux2_2
XFILLER_0_168_241 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14683_ VGND VPWR VGND VPWR _09137_ _09646_ _09036_ _09145_ _10150_ sky130_fd_sc_hd__o22a_2
XFILLER_0_135_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11895_ VGND VPWR result[114] _07511_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_39_420 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_196_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19210_ VPWR VGND keymem.key_mem\[13\]\[62\] _04972_ _04961_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16422_ VPWR VGND VGND VPWR _02580_ _02581_ _02582_ _02583_ _02584_ sky130_fd_sc_hd__and4b_2
XFILLER_0_32_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13634_ VGND VPWR _09106_ _09105_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_41_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_924 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_128_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_131_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16353_ VPWR VGND VGND VPWR _11308_ _02516_ _11316_ sky130_fd_sc_hd__nor2_2
XFILLER_0_27_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19141_ VGND VPWR VPWR VGND _04928_ _04927_ keymem.key_mem\[13\]\[36\] _04929_ sky130_fd_sc_hd__mux2_2
X_13565_ VGND VPWR VGND VPWR _09029_ _09016_ _09036_ _09033_ _09037_ sky130_fd_sc_hd__o22a_2
XFILLER_0_211_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15304_ VGND VPWR VGND VPWR _10766_ _10765_ _10764_ _10536_ sky130_fd_sc_hd__and3b_2
X_12516_ VPWR VGND VPWR VGND _08082_ keymem.key_mem\[10\]\[36\] _07629_ keymem.key_mem\[1\]\[36\]
+ _07969_ _08083_ sky130_fd_sc_hd__a221o_2
X_19072_ VPWR VGND keymem.key_mem_we _04889_ _10369_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16284_ VGND VPWR VGND VPWR _11211_ _11376_ _11527_ _11422_ _11323_ _02448_ sky130_fd_sc_hd__o32a_2
XFILLER_0_246_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_164_1200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13496_ VPWR VGND VPWR VGND _08968_ enc_block.block_w0_reg\[1\] _08952_ sky130_fd_sc_hd__or2_2
XFILLER_0_124_322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_48_1027 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15235_ VPWR VGND VGND VPWR _10595_ _10698_ _10516_ sky130_fd_sc_hd__nor2_2
X_18023_ VGND VPWR VGND VPWR _00272_ _03946_ _03945_ enc_block.round\[3\] sky130_fd_sc_hd__o21a_2
XFILLER_0_48_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12447_ VGND VPWR _08020_ _07662_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_50_640 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_23_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15166_ VGND VPWR VGND VPWR _10455_ _10575_ _10629_ _10490_ _10630_ sky130_fd_sc_hd__o22a_2
X_12378_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[24\] _07695_ keymem.key_mem\[9\]\[24\]
+ _07919_ _07957_ sky130_fd_sc_hd__a22o_2
XFILLER_0_151_196 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_142_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_386 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14117_ VPWR VGND VPWR VGND _09578_ _09587_ _09584_ _09575_ _09588_ sky130_fd_sc_hd__or4_2
XFILLER_0_1_269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15097_ VPWR VGND VGND VPWR _10561_ _10555_ _10560_ sky130_fd_sc_hd__nand2_2
XFILLER_0_103_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19974_ VPWR VGND VGND VPWR _05403_ keymem.key_mem\[10\]\[11\] _05402_ sky130_fd_sc_hd__nand2_2
XFILLER_0_205_1285 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_142_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_226_407 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18925_ VGND VPWR _04763_ enc_block.block_w0_reg\[10\] _04762_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_14048_ VGND VPWR _09520_ keymem.prev_key1_reg\[0\] keymem.prev_key1_reg\[32\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18856_ VGND VPWR _04701_ enc_block.block_w0_reg\[10\] enc_block.block_w0_reg\[15\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17807_ VPWR VGND VPWR VGND _03159_ _03800_ keymem.prev_key0_reg\[61\] _03788_ _00202_
+ sky130_fd_sc_hd__a22o_2
X_18787_ VGND VPWR _04639_ _04637_ _04638_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15999_ VGND VPWR _11454_ keymem.prev_key1_reg\[17\] keymem.prev_key1_reg\[49\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_253_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17738_ VGND VPWR VPWR VGND _03719_ key[164] keymem.prev_key1_reg\[36\] _03757_ sky130_fd_sc_hd__mux2_2
XFILLER_0_106_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17669_ VGND VPWR VPWR VGND _03691_ key[143] keymem.prev_key1_reg\[15\] _03709_ sky130_fd_sc_hd__mux2_2
X_19408_ VPWR VGND keymem.key_mem\[12\]\[4\] _05100_ _05095_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_15_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_127_1_Right_728 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20680_ VGND VPWR _01100_ _05775_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_110_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_358 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1042 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19339_ VGND VPWR _00481_ _05053_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_905 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_174_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_72_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22350_ VGND VPWR _01880_ _06665_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_169_1188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_286 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21301_ VGND VPWR VPWR VGND _06098_ _03633_ keymem.key_mem\[6\]\[122\] _06107_ sky130_fd_sc_hd__mux2_2
XFILLER_0_142_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22281_ VGND VPWR _01847_ _06629_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_13_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_115_388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_597 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24020_ VGND VPWR VPWR VGND clk _00513_ reset_n keymem.key_mem\[12\]\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_130_325 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21232_ VGND VPWR VPWR VGND _06065_ _03409_ keymem.key_mem\[6\]\[89\] _06071_ sky130_fd_sc_hd__mux2_2
XFILLER_0_198_76 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_130_336 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21163_ VGND VPWR VPWR VGND _06029_ _03108_ keymem.key_mem\[6\]\[56\] _06035_ sky130_fd_sc_hd__mux2_2
XFILLER_0_106_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20114_ VGND VPWR VPWR VGND _05469_ _03314_ keymem.key_mem\[10\]\[78\] _05476_ sky130_fd_sc_hd__mux2_2
X_21094_ VGND VPWR VPWR VGND _05996_ _02660_ keymem.key_mem\[6\]\[23\] _05999_ sky130_fd_sc_hd__mux2_2
X_20045_ VGND VPWR VPWR VGND _05435_ _03006_ keymem.key_mem\[10\]\[45\] _05440_ sky130_fd_sc_hd__mux2_2
X_24922_ VGND VPWR VPWR VGND clk _01415_ reset_n keymem.key_mem\[5\]\[19\] sky130_fd_sc_hd__dfrtp_2
X_24853_ VGND VPWR VPWR VGND clk _01346_ reset_n keymem.key_mem\[6\]\[78\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_99_139 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_77_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23804_ VGND VPWR VPWR VGND clk _00297_ reset_n enc_block.block_w0_reg\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_198_859 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_213_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24784_ VGND VPWR VPWR VGND clk _01277_ reset_n keymem.key_mem\[6\]\[9\] sky130_fd_sc_hd__dfrtp_2
X_21996_ VGND VPWR VGND VPWR _06478_ keymem.key_mem_we _03162_ _06475_ _01713_ sky130_fd_sc_hd__a31o_2
XFILLER_0_241_999 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_233_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_318 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23735_ keymem.prev_key0_reg\[91\] clk _00232_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20947_ VGND VPWR VGND VPWR _05920_ keymem.key_mem_we _03347_ _05916_ _01222_ sky130_fd_sc_hd__a31o_2
XFILLER_0_221_690 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11680_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[7\] dec_new_block\[7\]
+ _07404_ sky130_fd_sc_hd__mux2_2
X_23666_ keymem.prev_key0_reg\[22\] clk _00163_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20878_ VGND VPWR _01190_ _05883_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_165_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_95_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_187_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25405_ VGND VPWR VPWR VGND clk _01898_ reset_n keymem.key_mem\[2\]\[118\] sky130_fd_sc_hd__dfrtp_2
X_22617_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[127\] _06756_ _03793_ _05089_ _02035_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_14_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23597_ VGND VPWR VPWR VGND clk _00098_ reset_n keymem.key_mem\[14\]\[86\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_180_214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25336_ VGND VPWR VPWR VGND clk _01829_ reset_n keymem.key_mem\[2\]\[49\] sky130_fd_sc_hd__dfrtp_2
X_13350_ VPWR VGND VPWR VGND _08834_ keymem.key_mem\[6\]\[118\] _07657_ keymem.key_mem\[10\]\[118\]
+ _07909_ _08835_ sky130_fd_sc_hd__a221o_2
XFILLER_0_187_1277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22548_ VPWR VGND VGND VPWR _06761_ keymem.key_mem\[1\]\[75\] _06756_ sky130_fd_sc_hd__nand2_2
XFILLER_0_148_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_247 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_84_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12301_ VPWR VGND VPWR VGND _07885_ keymem.key_mem\[5\]\[18\] _07613_ keymem.key_mem\[9\]\[18\]
+ _07612_ _07886_ sky130_fd_sc_hd__a221o_2
X_13281_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[111\] _07597_ keymem.key_mem\[1\]\[111\]
+ _07969_ _08773_ sky130_fd_sc_hd__a22o_2
X_25267_ VGND VPWR VPWR VGND clk _01760_ reset_n keymem.key_mem\[3\]\[108\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22479_ VGND VPWR VPWR VGND _06726_ keymem.key_mem\[1\]\[34\] _02894_ _06733_ sky130_fd_sc_hd__mux2_2
XFILLER_0_32_640 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15020_ VPWR VGND VPWR VGND _10483_ _10464_ _10463_ _10472_ _10484_ sky130_fd_sc_hd__or4_2
XFILLER_0_32_651 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24218_ VGND VPWR VPWR VGND clk _00711_ reset_n keymem.key_mem\[11\]\[83\] sky130_fd_sc_hd__dfrtp_2
X_12232_ VGND VPWR enc_block.round_key\[12\] _07822_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_224_1149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25198_ VGND VPWR VPWR VGND clk _01691_ reset_n keymem.key_mem\[3\]\[39\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_993 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24149_ VGND VPWR VPWR VGND clk _00642_ reset_n keymem.key_mem\[11\]\[14\] sky130_fd_sc_hd__dfrtp_2
X_12163_ VPWR VGND VPWR VGND _07757_ keymem.key_mem\[13\]\[8\] _07588_ keymem.key_mem\[10\]\[8\]
+ _07562_ _07758_ sky130_fd_sc_hd__a221o_2
XFILLER_0_31_194 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_124_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16971_ VGND VPWR VPWR VGND _03084_ keymem.key_mem\[14\]\[55\] _03099_ _03100_ sky130_fd_sc_hd__mux2_2
X_12094_ VGND VPWR _07692_ _07550_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18710_ VGND VPWR _04569_ enc_block.block_w0_reg\[5\] _04363_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_159_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15922_ VGND VPWR VPWR VGND _11377_ _11345_ _11376_ _11378_ sky130_fd_sc_hd__or3_2
X_19690_ VGND VPWR VPWR VGND _05247_ keymem.key_mem\[11\]\[6\] _10284_ _05252_ sky130_fd_sc_hd__mux2_2
XFILLER_0_36_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1259 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18641_ VGND VPWR _04508_ _04373_ _04507_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15853_ VGND VPWR VGND VPWR _11245_ _11303_ _11308_ _11306_ _11309_ sky130_fd_sc_hd__o22a_2
XFILLER_0_95_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1223 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_243_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_239_1392 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_56_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_955 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14804_ VGND VPWR VGND VPWR _09517_ _10268_ _10266_ _10267_ _10270_ sky130_fd_sc_hd__a31o_2
XFILLER_0_235_1245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18572_ VPWR VGND VPWR VGND _04446_ _04443_ _04445_ sky130_fd_sc_hd__or2_2
X_15784_ VGND VPWR VPWR VGND _11173_ _11216_ _11233_ _11240_ sky130_fd_sc_hd__or3_2
X_12996_ VPWR VGND VPWR VGND _08515_ keymem.key_mem\[7\]\[83\] _07609_ keymem.key_mem\[10\]\[83\]
+ _07865_ _08516_ sky130_fd_sc_hd__a221o_2
XFILLER_0_54_1020 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_515 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_54_1031 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17523_ VPWR VGND _09533_ _03591_ _03590_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_8_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14735_ VGND VPWR VGND VPWR _09675_ _10169_ _10201_ _10200_ _09936_ sky130_fd_sc_hd__nor4_2
X_11947_ VGND VPWR _07550_ _07549_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14666_ VPWR VGND VGND VPWR _09420_ _09754_ _09441_ _09466_ _10133_ _10132_ sky130_fd_sc_hd__o221a_2
X_17454_ VPWR VGND VGND VPWR _03531_ _03532_ keylen sky130_fd_sc_hd__nor2_2
X_11878_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[10\] dec_new_block\[106\]
+ _07503_ sky130_fd_sc_hd__mux2_2
X_16405_ VGND VPWR VGND VPWR _11239_ _11466_ _11332_ _11400_ _02567_ sky130_fd_sc_hd__o22a_2
X_13617_ VGND VPWR _09089_ _09088_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14597_ VPWR VGND VPWR VGND _10062_ _10064_ _10063_ _09325_ _10065_ sky130_fd_sc_hd__or4_2
X_17385_ VGND VPWR VPWR VGND _09927_ _03471_ key[225] _03472_ sky130_fd_sc_hd__mux2_2
XFILLER_0_229_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19124_ VPWR VGND keymem.key_mem\[13\]\[30\] _04918_ _04915_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16336_ VGND VPWR VGND VPWR _02455_ _11377_ _11291_ _11357_ _02499_ sky130_fd_sc_hd__a31o_2
XFILLER_0_54_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13548_ VPWR VGND VGND VPWR _09019_ _09020_ _09016_ sky130_fd_sc_hd__nor2_2
XFILLER_0_166_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16267_ VPWR VGND VGND VPWR _11316_ _11204_ _02431_ _11399_ _11282_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_124_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19055_ VGND VPWR VPWR VGND keymem.round_ctr_reg\[1\] _09538_ _07387_ _04879_ sky130_fd_sc_hd__or3_2
XFILLER_0_2_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13479_ VPWR VGND VPWR VGND _08951_ enc_block.sword_ctr_reg\[0\] enc_block.sword_ctr_reg\[1\]
+ sky130_fd_sc_hd__or2_2
XFILLER_0_242_1205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15218_ VPWR VGND VPWR VGND _10499_ _10678_ _10679_ _10680_ _10681_ sky130_fd_sc_hd__or4bb_2
X_18006_ VGND VPWR VGND VPWR _03936_ _03935_ _03675_ _03652_ sky130_fd_sc_hd__and3b_2
XFILLER_0_23_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16198_ VPWR VGND VPWR VGND _02358_ _02362_ _02361_ _02356_ _02363_ sky130_fd_sc_hd__or4_2
XFILLER_0_112_358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_267_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15149_ VGND VPWR VGND VPWR _10608_ _10609_ _10522_ _10612_ _10613_ sky130_fd_sc_hd__o22a_2
XFILLER_0_205_1060 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_103_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19957_ VGND VPWR _00759_ _05393_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_10_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18908_ VPWR VGND VPWR VGND _04748_ _04684_ _04746_ sky130_fd_sc_hd__or2_2
XFILLER_0_177_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19888_ VGND VPWR _00728_ _05355_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_78_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_177_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18839_ VGND VPWR _04686_ _04683_ _04685_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21850_ VGND VPWR _01648_ _06397_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_218_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20801_ VPWR VGND keymem.key_mem\[7\]\[15\] _05842_ _05830_ VPWR VGND sky130_fd_sc_hd__and2_2
X_21781_ VGND VPWR _01615_ _06361_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_222_498 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23520_ VGND VPWR VPWR VGND clk _00021_ reset_n keymem.key_mem\[14\]\[9\] sky130_fd_sc_hd__dfrtp_2
X_20732_ VGND VPWR _01125_ _05802_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_92_304 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_77_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_100_1_Left_367 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_114_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_412 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_188_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23451_ VPWR VGND VGND VPWR _07192_ _07317_ _04248_ sky130_fd_sc_hd__nor2_2
XFILLER_0_11_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_128_1_Right_729 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20663_ VGND VPWR _01092_ _05766_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_149_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_188_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22402_ VGND VPWR _01905_ _06692_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_34_916 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_85_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23382_ VPWR VGND VPWR VGND _07255_ _04874_ _07254_ enc_block.block_w3_reg\[17\]
+ _07115_ _02322_ sky130_fd_sc_hd__a221o_2
XFILLER_0_184_1428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_489 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20594_ VGND VPWR _01059_ _05730_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_149_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25121_ VGND VPWR VPWR VGND clk _01614_ reset_n keymem.key_mem\[4\]\[90\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_229_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_85_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22333_ VGND VPWR _01872_ _06656_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_46_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_264_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25052_ VGND VPWR VPWR VGND clk _01545_ reset_n keymem.key_mem\[4\]\[21\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22264_ VGND VPWR _01839_ _06620_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_44_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_225_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24003_ VGND VPWR VPWR VGND clk _00496_ reset_n keymem.key_mem\[13\]\[124\] sky130_fd_sc_hd__dfrtp_2
X_21215_ VGND VPWR VPWR VGND _06052_ _03339_ keymem.key_mem\[6\]\[81\] _06062_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_130_2_Left_601 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22195_ VGND VPWR _01806_ _06584_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_223_1171 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_121_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21146_ VGND VPWR VPWR VGND _06018_ _03035_ keymem.key_mem\[6\]\[48\] _06026_ sky130_fd_sc_hd__mux2_2
XFILLER_0_79_1307 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_245_524 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21077_ VGND VPWR VPWR VGND _05983_ _11148_ keymem.key_mem\[6\]\[15\] _05990_ sky130_fd_sc_hd__mux2_2
XFILLER_0_156_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20028_ VGND VPWR VPWR VGND _05424_ _02924_ keymem.key_mem\[10\]\[37\] _05431_ sky130_fd_sc_hd__mux2_2
X_24905_ VGND VPWR VPWR VGND clk _01398_ reset_n keymem.key_mem\[5\]\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_236_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12850_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[68\] _08124_ _08384_ _08380_ _08385_
+ sky130_fd_sc_hd__o22a_2
X_24836_ VGND VPWR VPWR VGND clk _01329_ reset_n keymem.key_mem\[6\]\[61\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_236_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11801_ VGND VPWR result[67] _07464_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12781_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[61\] _07644_ _08322_ _08318_ _08323_
+ sky130_fd_sc_hd__o22a_2
X_24767_ VGND VPWR VPWR VGND clk _01260_ reset_n keymem.key_mem\[7\]\[120\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21979_ VGND VPWR _06469_ _06405_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_240_295 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_185_328 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14520_ VGND VPWR VGND VPWR _09985_ _09988_ _09989_ _09934_ sky130_fd_sc_hd__nand3_2
X_11732_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[1\] dec_new_block\[33\]
+ _07430_ sky130_fd_sc_hd__mux2_2
XFILLER_0_90_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23718_ keymem.prev_key0_reg\[74\] clk _00215_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_24698_ VGND VPWR VPWR VGND clk _01191_ reset_n keymem.key_mem\[7\]\[51\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_132_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14451_ VPWR VGND VGND VPWR _09576_ _09920_ _09358_ sky130_fd_sc_hd__nor2_2
X_23649_ keymem.prev_key0_reg\[5\] clk _00146_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_11663_ VPWR VGND VPWR VGND aes_core_ctrl_reg\[2\] _07371_ init aes_core_ctrl_reg\[0\]
+ _00006_ sky130_fd_sc_hd__a22o_2
XFILLER_0_3_1057 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13402_ VPWR VGND VPWR VGND _08881_ keymem.key_mem\[6\]\[123\] _07759_ keymem.key_mem\[8\]\[123\]
+ _07752_ _08882_ sky130_fd_sc_hd__a221o_2
XFILLER_0_193_383 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_125_2_Left_596 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17170_ VPWR VGND VGND VPWR _03280_ keymem.key_mem\[14\]\[74\] _09541_ sky130_fd_sc_hd__nand2_2
XFILLER_0_153_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14382_ VGND VPWR VGND VPWR _09789_ _09759_ keymem.round_ctr_reg\[0\] _09852_ sky130_fd_sc_hd__a21o_2
XFILLER_0_24_404 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_64_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16121_ VGND VPWR VGND VPWR _11296_ _11238_ _11352_ _11422_ _11323_ _11575_ sky130_fd_sc_hd__o32a_2
XFILLER_0_88_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25319_ VGND VPWR VPWR VGND clk _01812_ reset_n keymem.key_mem\[2\]\[32\] sky130_fd_sc_hd__dfrtp_2
X_13333_ VGND VPWR VGND VPWR _08096_ keymem.key_mem\[5\]\[116\] _08815_ _08817_ _08820_
+ _08819_ sky130_fd_sc_hd__a2111o_2
XPHY_EDGE_ROW_94_1_Left_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_49_1166 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_51_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_243_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16052_ VPWR VGND VPWR VGND _11506_ _11357_ _11348_ _11427_ _11434_ _11507_ sky130_fd_sc_hd__a221o_2
X_13264_ VPWR VGND VPWR VGND _08757_ keymem.key_mem\[11\]\[109\] _07838_ keymem.key_mem\[4\]\[109\]
+ _07552_ _08758_ sky130_fd_sc_hd__a221o_2
XFILLER_0_204_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15003_ VGND VPWR VPWR VGND _10453_ _10466_ _10451_ _10467_ sky130_fd_sc_hd__or3_2
XFILLER_0_267_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12215_ VGND VPWR _07806_ _07577_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_161_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13195_ VGND VPWR enc_block.round_key\[102\] _08695_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_202_1200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19811_ VGND VPWR _00691_ _05315_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12146_ VGND VPWR _07742_ _07560_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_102_391 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19742_ VGND VPWR VPWR VGND _05270_ keymem.key_mem\[11\]\[31\] _02862_ _05279_ sky130_fd_sc_hd__mux2_2
X_16954_ VGND VPWR VPWR VGND _03084_ keymem.key_mem\[14\]\[53\] _03083_ _03085_ sky130_fd_sc_hd__mux2_2
X_12077_ VGND VPWR VGND VPWR _07677_ _07665_ keymem.key_mem\[4\]\[3\] _07669_ _07676_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_47_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15905_ VGND VPWR _11361_ _11360_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19673_ keymem.round_ctr_reg\[0\] _05241_ keymem.key_mem_we keymem.round_ctr_reg\[1\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_16885_ VPWR VGND VPWR VGND _11110_ _03022_ _11144_ _11624_ sky130_fd_sc_hd__or3b_2
XFILLER_0_217_793 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_205_933 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_204_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18624_ VPWR VGND VPWR VGND _04492_ block[83] _04487_ enc_block.block_w2_reg\[19\]
+ _04425_ _04493_ sky130_fd_sc_hd__a221o_2
X_15836_ VGND VPWR VGND VPWR _11292_ _11229_ _11228_ _11272_ _11226_ sky130_fd_sc_hd__and4_2
XFILLER_0_59_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_59_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18555_ VPWR VGND VPWR VGND _04430_ block[76] _04330_ enc_block.block_w3_reg\[12\]
+ _04425_ _04431_ sky130_fd_sc_hd__a221o_2
XFILLER_0_188_166 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15767_ VPWR VGND VGND VPWR _11174_ _11223_ _11167_ sky130_fd_sc_hd__nor2_2
X_12979_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[81\] _07651_ keymem.key_mem\[1\]\[81\]
+ _07670_ _08501_ sky130_fd_sc_hd__a22o_2
XFILLER_0_176_317 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_172_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17506_ VPWR VGND _11553_ _03576_ _11554_ VPWR VGND sky130_fd_sc_hd__and2_2
X_14718_ VPWR VGND VGND VPWR _10185_ _10168_ _10184_ sky130_fd_sc_hd__nand2_2
X_18486_ VPWR VGND VPWR VGND _04368_ block[69] _04330_ enc_block.block_w0_reg\[5\]
+ _04276_ _04369_ sky130_fd_sc_hd__a221o_2
XFILLER_0_86_175 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15698_ VGND VPWR keymem.prev_key1_reg\[80\] _11152_ _11154_ _11153_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_170_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_86_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17437_ VPWR VGND VGND VPWR _03516_ _03517_ keylen sky130_fd_sc_hd__nor2_2
X_14649_ VGND VPWR VGND VPWR _09327_ _09323_ _09403_ _09495_ _10116_ sky130_fd_sc_hd__o22a_2
XFILLER_0_27_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_916 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_55_551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_129_299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_573 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17368_ VGND VPWR VGND VPWR _02855_ _02854_ _09866_ _03457_ sky130_fd_sc_hd__a21o_2
XFILLER_0_103_74 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_437 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19107_ VPWR VGND keymem.key_mem\[13\]\[22\] _04909_ _04903_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16319_ VPWR VGND VPWR VGND _02482_ keymem.prev_key1_reg\[21\] sky130_fd_sc_hd__inv_2
XFILLER_0_67_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17299_ VPWR VGND VPWR VGND _03395_ keymem.prev_key0_reg\[88\] sky130_fd_sc_hd__inv_2
XFILLER_0_28_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19038_ VPWR VGND VPWR VGND _04863_ _04505_ enc_block.block_w2_reg\[30\] _04504_
+ _04864_ sky130_fd_sc_hd__a22o_2
XFILLER_0_259_627 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_854 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_152_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1166 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_11_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21000_ VGND VPWR VPWR VGND _05945_ _05050_ keymem.key_mem\[7\]\[108\] _05948_ sky130_fd_sc_hd__mux2_2
XFILLER_0_10_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_255_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_49_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_214_218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22951_ VGND VPWR VGND VPWR _06938_ _02868_ _02865_ _02871_ _06892_ sky130_fd_sc_hd__a211o_2
XFILLER_0_138_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21902_ VPWR VGND keymem.key_mem\[3\]\[18\] _06428_ _06427_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_78_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1251 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25670_ VGND VPWR VPWR VGND clk _02163_ reset_n keymem.key_mem\[0\]\[127\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22882_ VGND VPWR VGND VPWR _10271_ _06890_ _10282_ _06895_ sky130_fd_sc_hd__a21o_2
XFILLER_0_223_763 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_190_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24621_ VGND VPWR VPWR VGND clk _01114_ reset_n keymem.key_mem\[8\]\[102\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_250_582 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21833_ VGND VPWR VPWR VGND _06388_ _03592_ keymem.key_mem\[4\]\[116\] _06389_ sky130_fd_sc_hd__mux2_2
XFILLER_0_190_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24552_ VGND VPWR VPWR VGND clk _01045_ reset_n keymem.key_mem\[8\]\[33\] sky130_fd_sc_hd__dfrtp_2
X_21764_ VGND VPWR _01607_ _06352_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23503_ VGND VPWR VGND VPWR _07361_ enc_block.round_key\[31\] _04148_ _07363_ sky130_fd_sc_hd__a21o_2
XFILLER_0_182_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_65_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20715_ VGND VPWR _01117_ _05793_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24483_ VGND VPWR VPWR VGND clk _00976_ reset_n keymem.key_mem\[9\]\[92\] sky130_fd_sc_hd__dfrtp_2
X_21695_ VGND VPWR _01574_ _06316_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_18_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23434_ VGND VPWR VGND VPWR _07302_ _04064_ _07301_ _07300_ sky130_fd_sc_hd__o21a_2
XFILLER_0_92_167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20646_ VGND VPWR _01084_ _05757_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_190_342 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_595 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23365_ VPWR VGND VPWR VGND _07240_ enc_block.block_w0_reg\[23\] _07239_ sky130_fd_sc_hd__or2_2
X_20577_ VGND VPWR _01051_ _05721_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_46_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1102 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25104_ VGND VPWR VPWR VGND clk _01597_ reset_n keymem.key_mem\[4\]\[73\] sky130_fd_sc_hd__dfrtp_2
X_22316_ VGND VPWR VPWR VGND _06647_ _03364_ keymem.key_mem\[2\]\[84\] _06648_ sky130_fd_sc_hd__mux2_2
X_23296_ VPWR VGND VGND VPWR _07177_ _07178_ _07175_ sky130_fd_sc_hd__nor2_2
XFILLER_0_14_470 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_239_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1266 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25035_ VGND VPWR VPWR VGND clk _01528_ reset_n keymem.key_mem\[4\]\[4\] sky130_fd_sc_hd__dfrtp_2
X_22247_ VGND VPWR VPWR VGND _06611_ _03067_ keymem.key_mem\[2\]\[51\] _06612_ sky130_fd_sc_hd__mux2_2
X_12000_ VGND VPWR _07603_ _07602_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22178_ VGND VPWR _01798_ _06575_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21129_ VGND VPWR VPWR VGND _06007_ _02955_ keymem.key_mem\[6\]\[40\] _06017_ sky130_fd_sc_hd__mux2_2
XFILLER_0_233_516 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13951_ VGND VPWR _09423_ _09422_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_96_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12902_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[74\] _07779_ keymem.key_mem\[14\]\[74\]
+ _08003_ _08431_ sky130_fd_sc_hd__a22o_2
X_13882_ VPWR VGND VPWR VGND _09307_ _09291_ _09285_ _09306_ _09354_ sky130_fd_sc_hd__or4_2
X_16670_ VGND VPWR _02824_ keymem.prev_key0_reg\[62\] keymem.prev_key0_reg\[94\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15621_ VGND VPWR VGND VPWR _11078_ _10718_ _11079_ _10580_ sky130_fd_sc_hd__a21oi_2
X_12833_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[67\] _07591_ keymem.key_mem\[2\]\[67\]
+ _07545_ _08369_ sky130_fd_sc_hd__a22o_2
X_24819_ VGND VPWR VPWR VGND clk _01312_ reset_n keymem.key_mem\[6\]\[44\] sky130_fd_sc_hd__dfrtp_2
X_25799_ keymem.prev_key1_reg\[115\] clk _02292_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_33_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18340_ VPWR VGND VPWR VGND _04237_ block[120] _04213_ enc_block.block_w0_reg\[24\]
+ _04171_ _04238_ sky130_fd_sc_hd__a221o_2
X_15552_ VPWR VGND VGND VPWR _10587_ _11011_ _10449_ sky130_fd_sc_hd__nor2_2
X_12764_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[60\] _07649_ keymem.key_mem\[4\]\[60\]
+ _07913_ _08307_ sky130_fd_sc_hd__a22o_2
XFILLER_0_51_1045 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_68_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_185_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_1056 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14503_ VGND VPWR VGND VPWR _09972_ _09971_ _09968_ _09967_ _09807_ sky130_fd_sc_hd__and4_2
XFILLER_0_68_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11715_ VGND VPWR result[24] _07421_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15483_ VGND VPWR VPWR VGND _10943_ _10475_ _10672_ _10541_ _10942_ sky130_fd_sc_hd__o31a_2
X_18271_ VPWR VGND VPWR VGND _04175_ _04089_ _04173_ sky130_fd_sc_hd__or2_2
X_12695_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[53\] _07668_ keymem.key_mem\[4\]\[53\]
+ _07734_ _08245_ sky130_fd_sc_hd__a22o_2
XFILLER_0_12_1029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17222_ VPWR VGND VPWR VGND _03326_ key[80] _08935_ sky130_fd_sc_hd__or2_2
X_14434_ VPWR VGND VGND VPWR _09431_ _09422_ _09903_ _09366_ _09418_ sky130_fd_sc_hd__o22ai_2
X_11646_ VPWR VGND VPWR VGND _00002_ _07383_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14365_ VGND VPWR VGND VPWR _09067_ _09178_ _09091_ _09148_ _09835_ sky130_fd_sc_hd__o22a_2
X_17153_ VPWR VGND VPWR VGND _03264_ key[73] _08935_ sky130_fd_sc_hd__or2_2
XFILLER_0_68_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_12_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16104_ VPWR VGND VPWR VGND _11558_ _11556_ _11557_ sky130_fd_sc_hd__or2_2
X_13316_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[115\] _08137_ keymem.key_mem\[10\]\[115\]
+ _07785_ _08804_ sky130_fd_sc_hd__a22o_2
X_17084_ VGND VPWR VPWR VGND _03185_ keymem.key_mem\[14\]\[65\] _03202_ _03203_ sky130_fd_sc_hd__mux2_2
XFILLER_0_208_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14296_ VPWR VGND VGND VPWR _09311_ _09353_ _09766_ _09386_ _09401_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_204_1317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_149_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16035_ VGND VPWR VPWR VGND _11485_ _11489_ _11481_ _11490_ sky130_fd_sc_hd__or3_2
X_13247_ VGND VPWR enc_block.round_key\[107\] _08742_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_208_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1163 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13178_ VPWR VGND VPWR VGND _08679_ keymem.key_mem\[10\]\[101\] _07909_ keymem.key_mem\[4\]\[101\]
+ _07914_ _08680_ sky130_fd_sc_hd__a221o_2
XFILLER_0_104_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12129_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[6\] _07674_ keymem.key_mem\[8\]\[6\]
+ _07540_ _07726_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_252_803 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17986_ VGND VPWR _00259_ _03922_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_263_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1096 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_139_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19725_ VGND VPWR _05270_ _05246_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_224_527 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16937_ VGND VPWR _00063_ _03069_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_139_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_346 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_252_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_261_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19656_ VGND VPWR VPWR VGND _05227_ _05075_ keymem.key_mem\[12\]\[120\] _05232_ sky130_fd_sc_hd__mux2_2
X_16868_ VGND VPWR VPWR VGND _02986_ keymem.key_mem\[14\]\[45\] _03006_ _03007_ sky130_fd_sc_hd__mux2_2
XFILLER_0_215_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18607_ VPWR VGND VPWR VGND _04477_ _04459_ _04476_ enc_block.block_w1_reg\[17\]
+ _04424_ _00325_ sky130_fd_sc_hd__a221o_2
XFILLER_0_204_262 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15819_ VPWR VGND VGND VPWR _11275_ _11167_ _11174_ sky130_fd_sc_hd__nand2_2
X_19587_ VPWR VGND keymem.key_mem\[12\]\[87\] _05196_ _05173_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_215_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16799_ VGND VPWR VGND VPWR _02941_ _10317_ _02942_ _02943_ _02944_ keylen sky130_fd_sc_hd__a221oi_2
XFILLER_0_149_328 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18538_ VPWR VGND VPWR VGND _04415_ _04291_ _04414_ enc_block.block_w1_reg\[10\]
+ _04317_ _00318_ sky130_fd_sc_hd__a221o_2
XFILLER_0_181_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_133_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_315 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_213_1170 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18469_ VGND VPWR _04353_ enc_block.block_w3_reg\[12\] _04352_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20500_ VGND VPWR _01014_ _05681_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_12_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21480_ VGND VPWR _01473_ _06202_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_16_724 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_56_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_146_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20431_ VGND VPWR VPWR VGND _05638_ _03485_ keymem.key_mem\[9\]\[99\] _05644_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_99_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_132_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23150_ VGND VPWR VGND VPWR _03552_ _03794_ _03554_ _07059_ sky130_fd_sc_hd__a21o_2
X_20362_ VGND VPWR VPWR VGND _05602_ _03209_ keymem.key_mem\[9\]\[66\] _05608_ sky130_fd_sc_hd__mux2_2
XFILLER_0_226_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22101_ VGND VPWR _01763_ _06533_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_3_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23081_ VGND VPWR VGND VPWR _07016_ _03361_ _06891_ _03363_ _07011_ sky130_fd_sc_hd__a211o_2
X_20293_ VGND VPWR VPWR VGND _05569_ _02883_ keymem.key_mem\[9\]\[33\] _05572_ sky130_fd_sc_hd__mux2_2
XFILLER_0_144_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22032_ VGND VPWR _01730_ _06497_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_11_473 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_215_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23983_ VGND VPWR VPWR VGND clk _00476_ reset_n keymem.key_mem\[13\]\[104\] sky130_fd_sc_hd__dfrtp_2
X_25722_ keymem.prev_key1_reg\[38\] clk _02215_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22934_ VGND VPWR VPWR VGND _02202_ _02707_ _02719_ _06925_ _06927_ sky130_fd_sc_hd__o31a_2
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_97_248 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22865_ VPWR VGND VPWR VGND _06883_ _09543_ _03672_ sky130_fd_sc_hd__or2_2
X_25653_ VGND VPWR VPWR VGND clk _02146_ reset_n keymem.key_mem\[0\]\[110\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_151_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24604_ VGND VPWR VPWR VGND clk _01097_ reset_n keymem.key_mem\[8\]\[85\] sky130_fd_sc_hd__dfrtp_2
X_21816_ VGND VPWR VPWR VGND _06377_ _03543_ keymem.key_mem\[4\]\[108\] _06380_ sky130_fd_sc_hd__mux2_2
XFILLER_0_190_1295 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25584_ VGND VPWR VPWR VGND clk _02077_ reset_n keymem.key_mem\[0\]\[41\] sky130_fd_sc_hd__dfrtp_2
X_22796_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[99\] _06850_ _06849_ _05031_ _02135_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_112_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_151_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24535_ VGND VPWR VPWR VGND clk _01028_ reset_n keymem.key_mem\[8\]\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_241_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21747_ VGND VPWR VGND VPWR _06259_ _03286_ _01599_ _06343_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_4_1141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_307 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12480_ VGND VPWR _08050_ _07748_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24466_ VGND VPWR VPWR VGND clk _00959_ reset_n keymem.key_mem\[9\]\[75\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21678_ VGND VPWR _01566_ _06307_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23417_ _07285_ _07287_ _04064_ _07286_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_20629_ VGND VPWR VPWR VGND _05747_ _03193_ keymem.key_mem\[8\]\[64\] _05749_ sky130_fd_sc_hd__mux2_2
XFILLER_0_123_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24397_ VGND VPWR VPWR VGND clk _00890_ reset_n keymem.key_mem\[9\]\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_163_386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14150_ VGND VPWR VGND VPWR _09621_ _09464_ _09371_ _09489_ _09370_ sky130_fd_sc_hd__and4_2
X_23348_ VPWR VGND VPWR VGND _07225_ _07148_ _07223_ sky130_fd_sc_hd__or2_2
XFILLER_0_22_749 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_162_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13101_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[93\] _07694_ keymem.key_mem\[1\]\[93\]
+ _07670_ _08611_ sky130_fd_sc_hd__a22o_2
XFILLER_0_0_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14081_ VPWR VGND VGND VPWR _09552_ _09361_ _09247_ sky130_fd_sc_hd__nand2_2
X_23279_ VPWR VGND VPWR VGND _07162_ block[7] _04837_ enc_block.block_w2_reg\[7\]
+ _04798_ _07163_ sky130_fd_sc_hd__a221o_2
XFILLER_0_162_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13032_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[86\] _08449_ _08548_ _08544_ _08549_
+ sky130_fd_sc_hd__o22a_2
X_25018_ VGND VPWR VPWR VGND clk _01511_ reset_n keymem.key_mem\[5\]\[115\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_30_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_265_438 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17840_ VGND VPWR VPWR VGND _03812_ key[200] keymem.prev_key1_reg\[72\] _03823_ sky130_fd_sc_hd__mux2_2
XFILLER_0_218_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_696 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17771_ VGND VPWR _00190_ _03776_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14983_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[8\] _10402_ _10447_ _09255_ _10395_
+ _10396_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_260_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_261_644 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19510_ VPWR VGND keymem.key_mem\[12\]\[51\] _05155_ _05128_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_260_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16722_ VGND VPWR VPWR VGND _02662_ keymem.key_mem\[14\]\[32\] _02873_ _02874_ sky130_fd_sc_hd__mux2_2
X_13934_ VPWR VGND VGND VPWR _09396_ _09397_ _09378_ _09330_ _09406_ _09405_ sky130_fd_sc_hd__o221a_2
XFILLER_0_44_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19441_ VPWR VGND keymem.key_mem\[12\]\[19\] _05118_ _05116_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_173_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16653_ VPWR VGND VGND VPWR _09732_ _02808_ key[157] sky130_fd_sc_hd__nor2_2
X_13865_ VGND VPWR VGND VPWR _09337_ _09274_ _09272_ keymem.prev_key1_reg\[31\] _08955_
+ _08942_ sky130_fd_sc_hd__a32o_2
X_15604_ VGND VPWR VPWR VGND _11060_ _11061_ _11059_ _11062_ sky130_fd_sc_hd__or3_2
X_12816_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[65\] _07924_ keymem.key_mem\[2\]\[65\]
+ _08131_ _08354_ sky130_fd_sc_hd__a22o_2
X_19372_ VGND VPWR VPWR VGND _05067_ _05075_ keymem.key_mem\[13\]\[120\] _05076_ sky130_fd_sc_hd__mux2_2
XFILLER_0_201_254 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16584_ VPWR VGND VPWR VGND _02741_ _02677_ _02732_ key[154] _02723_ _02742_ sky130_fd_sc_hd__a221o_2
X_13796_ VGND VPWR _09268_ _09267_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_70_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_130_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18323_ VGND VPWR VGND VPWR _02586_ _02572_ _04073_ _04223_ sky130_fd_sc_hd__a21o_2
XFILLER_0_134_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15535_ VGND VPWR _10580_ _10925_ _10994_ _10803_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_151_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_57_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12747_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[58\] _07838_ keymem.key_mem\[2\]\[58\]
+ _07816_ _08292_ sky130_fd_sc_hd__a22o_2
XFILLER_0_70_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18254_ VPWR VGND VGND VPWR _04159_ _04160_ _04041_ sky130_fd_sc_hd__nor2_2
X_15466_ VPWR VGND VGND VPWR _10627_ _10926_ _10522_ sky130_fd_sc_hd__nor2_2
XFILLER_0_44_329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12678_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[51\] _08145_ _08229_ _08225_ _08230_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_25_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17205_ VGND VPWR _02866_ key[78] _03311_ _03029_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_14417_ VPWR VGND VGND VPWR _09487_ _09886_ _09336_ sky130_fd_sc_hd__nor2_2
X_11629_ VGND VPWR aes_core_ctrl_reg\[0\] init _07370_ next VPWR VGND sky130_fd_sc_hd__o21ai_2
X_18185_ VPWR VGND VPWR VGND _04096_ _04040_ _04094_ enc_block.block_w0_reg\[10\]
+ _03976_ _00284_ sky130_fd_sc_hd__a221o_2
XFILLER_0_53_852 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15397_ VPWR VGND VGND VPWR _10629_ _10858_ _10511_ sky130_fd_sc_hd__nor2_2
XFILLER_0_29_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_180_1_Right_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_107_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17136_ VGND VPWR VGND VPWR _03249_ _09721_ _10732_ key[71] sky130_fd_sc_hd__o21a_2
X_14348_ VPWR VGND VGND VPWR _09103_ _09100_ _09110_ _09108_ _09818_ _09817_ sky130_fd_sc_hd__o221a_2
XFILLER_0_29_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_226 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_180_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_546 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_208_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14279_ VGND VPWR _09749_ _09623_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17067_ VPWR VGND VGND VPWR _03187_ key[192] _09522_ sky130_fd_sc_hd__nand2_2
XFILLER_0_141_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_180_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16018_ VGND VPWR _11473_ _11318_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_81_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_141_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_225_814 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_139_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_174_1202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_58_1018 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17969_ VGND VPWR VPWR VGND _03896_ _03910_ keymem.prev_key0_reg\[113\] _03911_ sky130_fd_sc_hd__mux2_2
X_19708_ VGND VPWR _00642_ _05261_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20980_ VGND VPWR _01238_ _05937_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_250_1101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19639_ VGND VPWR VPWR VGND _05216_ _05058_ keymem.key_mem\[12\]\[112\] _05223_ sky130_fd_sc_hd__mux2_2
XFILLER_0_191_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_149_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22650_ VGND VPWR VPWR VGND _06785_ keymem.key_mem\[0\]\[14\] _11099_ _06796_ sky130_fd_sc_hd__mux2_2
XFILLER_0_152_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_125_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21601_ VGND VPWR _01529_ _06267_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_149_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_657 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22581_ VGND VPWR _02003_ _06773_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24320_ VGND VPWR VPWR VGND clk _00813_ reset_n keymem.key_mem\[10\]\[57\] sky130_fd_sc_hd__dfrtp_2
X_21532_ VGND VPWR _01498_ _06229_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_1_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_185_1320 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_141_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1052 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24251_ VGND VPWR VPWR VGND clk _00744_ reset_n keymem.key_mem\[11\]\[116\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21463_ VGND VPWR _01465_ _06193_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_141_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23202_ VGND VPWR _07093_ _07092_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20414_ VGND VPWR VPWR VGND _05627_ _03427_ keymem.key_mem\[9\]\[91\] _05635_ sky130_fd_sc_hd__mux2_2
XFILLER_0_160_345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24182_ VGND VPWR VPWR VGND clk _00675_ reset_n keymem.key_mem\[11\]\[47\] sky130_fd_sc_hd__dfrtp_2
X_21394_ VGND VPWR _01432_ _06157_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_120_209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23133_ VGND VPWR _02281_ _07047_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_113_250 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20345_ VGND VPWR VPWR VGND _05591_ _03130_ keymem.key_mem\[9\]\[58\] _05599_ sky130_fd_sc_hd__mux2_2
XFILLER_0_222_1225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_1000 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23064_ VGND VPWR VGND VPWR _02254_ _07005_ _06954_ keymem.prev_key1_reg\[77\] sky130_fd_sc_hd__o21a_2
X_20276_ VGND VPWR VPWR VGND _05558_ _02721_ keymem.key_mem\[9\]\[25\] _05563_ sky130_fd_sc_hd__mux2_2
X_22015_ VGND VPWR _01722_ _06488_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_192_1335 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_58_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11980_ VGND VPWR _07583_ _07582_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23966_ VGND VPWR VPWR VGND clk _00459_ reset_n keymem.key_mem\[13\]\[87\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25705_ keymem.prev_key1_reg\[21\] clk _02198_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22917_ VGND VPWR _06916_ _06881_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23897_ VGND VPWR VPWR VGND clk _00390_ reset_n keymem.key_mem\[13\]\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_252_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_2_Left_542 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13650_ VGND VPWR _09122_ _09121_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25636_ VGND VPWR VPWR VGND clk _02129_ reset_n keymem.key_mem\[0\]\[93\] sky130_fd_sc_hd__dfrtp_2
X_22848_ VGND VPWR VGND VPWR _06872_ _06871_ _05530_ keymem.round_ctr_rst sky130_fd_sc_hd__and3b_2
XFILLER_0_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12601_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[44\] _07694_ keymem.key_mem\[12\]\[44\]
+ _07806_ _08160_ sky130_fd_sc_hd__a22o_2
XFILLER_0_13_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13581_ VGND VPWR _09053_ _09052_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_39_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22779_ VGND VPWR _02123_ _06851_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25567_ VGND VPWR VPWR VGND clk _02060_ reset_n keymem.key_mem\[0\]\[24\] sky130_fd_sc_hd__dfrtp_2
X_15320_ VPWR VGND VGND VPWR _10588_ _10782_ _10608_ sky130_fd_sc_hd__nor2_2
X_12532_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[38\] _08009_ keymem.key_mem\[6\]\[38\]
+ _07711_ _08097_ sky130_fd_sc_hd__a22o_2
XFILLER_0_13_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24518_ VGND VPWR VPWR VGND clk _01011_ reset_n keymem.key_mem\[9\]\[127\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26_329 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25498_ VGND VPWR VPWR VGND clk _01991_ reset_n keymem.key_mem\[1\]\[83\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15251_ VGND VPWR VPWR VGND _10478_ _10588_ _10580_ _10714_ sky130_fd_sc_hd__or3_2
X_12463_ VPWR VGND VPWR VGND _08034_ keymem.key_mem\[7\]\[31\] _07609_ keymem.key_mem\[9\]\[31\]
+ _07738_ _08035_ sky130_fd_sc_hd__a221o_2
XFILLER_0_163_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24449_ VGND VPWR VPWR VGND clk _00942_ reset_n keymem.key_mem\[9\]\[58\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_129_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14202_ VPWR VGND VGND VPWR _09132_ _09673_ _09174_ sky130_fd_sc_hd__nor2_2
X_15182_ VGND VPWR _10646_ _10465_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_22_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_919 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12394_ VPWR VGND VPWR VGND _07971_ keymem.key_mem\[6\]\[25\] _07711_ keymem.key_mem\[10\]\[25\]
+ _07743_ _07972_ sky130_fd_sc_hd__a221o_2
XFILLER_0_62_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_151_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14133_ VPWR VGND VGND VPWR _09301_ _09565_ _09604_ _09349_ _09486_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_209_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19990_ VGND VPWR VPWR VGND _05400_ _02410_ keymem.key_mem\[10\]\[19\] _05411_ sky130_fd_sc_hd__mux2_2
XFILLER_0_205_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_579 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18941_ VGND VPWR _04778_ _04599_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14064_ VGND VPWR VGND VPWR _08930_ key[128] _09535_ _09536_ sky130_fd_sc_hd__a21o_2
XFILLER_0_162_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13015_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[85\] _07787_ keymem.key_mem\[1\]\[85\]
+ _07714_ _08533_ sky130_fd_sc_hd__a22o_2
X_18872_ VPWR VGND _04716_ _04715_ enc_block.round_key\[44\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_20_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1268 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_158_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17823_ VGND VPWR VPWR VGND _03777_ _03810_ keymem.prev_key0_reg\[67\] _03811_ sky130_fd_sc_hd__mux2_2
XFILLER_0_94_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17754_ VGND VPWR VPWR VGND _03763_ _03766_ keymem.prev_key0_reg\[42\] _03767_ sky130_fd_sc_hd__mux2_2
X_14966_ VGND VPWR _10430_ _10429_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_55_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16705_ VGND VPWR VGND VPWR _02855_ _02854_ _02858_ _02856_ sky130_fd_sc_hd__a21oi_2
X_13917_ VGND VPWR VPWR VGND _09331_ _09246_ _09303_ _09389_ sky130_fd_sc_hd__or3_2
X_17685_ VGND VPWR VPWR VGND _03719_ key[148] keymem.prev_key1_reg\[20\] _03720_ sky130_fd_sc_hd__mux2_2
XFILLER_0_216_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14897_ VGND VPWR VGND VPWR _10315_ _10292_ keymem.round_ctr_reg\[0\] _10362_ sky130_fd_sc_hd__a21o_2
X_19424_ VGND VPWR _00511_ _05108_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_173_1290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16636_ _10108_ _02791_ keymem.round_ctr_reg\[0\] _10140_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_76_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13848_ VGND VPWR VGND VPWR _09320_ _09246_ _09300_ _09319_ _09304_ sky130_fd_sc_hd__a211o_2
XFILLER_0_134_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19355_ VPWR VGND keymem.key_mem_we _05064_ _03585_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_31_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16567_ VGND VPWR VGND VPWR _11618_ keymem.rcon_reg\[2\] _02725_ _11589_ sky130_fd_sc_hd__nand3_2
X_13779_ VGND VPWR VGND VPWR enc_block.block_w1_reg\[27\] _08985_ _09249_ _09022_
+ _09251_ _09250_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_35_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18306_ VGND VPWR VGND VPWR _04205_ _04204_ _04207_ _04203_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_224_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15518_ VGND VPWR VPWR VGND _09864_ keymem.key_mem\[14\]\[12\] _10977_ _10978_ sky130_fd_sc_hd__mux2_2
XFILLER_0_139_191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19286_ VGND VPWR VGND VPWR _05018_ keymem.key_mem_we _03427_ _04999_ _00463_ sky130_fd_sc_hd__a31o_2
X_16498_ VPWR VGND VPWR VGND _02656_ _02650_ _02659_ _02658_ keylen sky130_fd_sc_hd__a211oi_2
XFILLER_0_169_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_112_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18237_ VPWR VGND VPWR VGND _04144_ _04140_ _04142_ sky130_fd_sc_hd__or2_2
XFILLER_0_127_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15449_ VGND VPWR VPWR VGND _09729_ _10909_ key[139] _10910_ sky130_fd_sc_hd__mux2_2
XFILLER_0_26_863 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18168_ VGND VPWR _04081_ _04078_ _04080_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_384 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_245_1269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_181_1_Right_782 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_74 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1033 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17119_ VGND VPWR VGND VPWR _08930_ key[197] _03233_ _03234_ sky130_fd_sc_hd__a21o_2
XFILLER_0_142_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18099_ VPWR VGND _04018_ _04017_ enc_block.round_key\[99\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_40_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_96_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_229_416 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20130_ VGND VPWR _00841_ _05484_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_141_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_78 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20061_ VGND VPWR _00808_ _05448_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_29_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23820_ VGND VPWR VPWR VGND clk _00313_ reset_n enc_block.block_w1_reg\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_225_688 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23751_ keymem.prev_key0_reg\[107\] clk _00248_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20963_ VGND VPWR VGND VPWR _05928_ keymem.key_mem_we _03418_ _05916_ _01230_ sky130_fd_sc_hd__a31o_2
XFILLER_0_221_850 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22702_ VGND VPWR _06819_ _03864_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23682_ keymem.prev_key0_reg\[38\] clk _00179_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_113_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20894_ VPWR VGND keymem.key_mem\[7\]\[58\] _05892_ _05886_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_152_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25421_ VGND VPWR VPWR VGND clk _01914_ reset_n keymem.key_mem\[1\]\[6\] sky130_fd_sc_hd__dfrtp_2
X_22633_ VGND VPWR _02041_ _06787_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_113_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_402 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25352_ VGND VPWR VPWR VGND clk _01845_ reset_n keymem.key_mem\[2\]\[65\] sky130_fd_sc_hd__dfrtp_2
X_22564_ VGND VPWR _06766_ _03859_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_152_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_14_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_187_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21515_ VGND VPWR VPWR VGND _06220_ _03452_ keymem.key_mem\[5\]\[94\] _06221_ sky130_fd_sc_hd__mux2_2
X_24303_ VGND VPWR VPWR VGND clk _00796_ reset_n keymem.key_mem\[10\]\[40\] sky130_fd_sc_hd__dfrtp_2
X_25283_ VGND VPWR VPWR VGND clk _01776_ reset_n keymem.key_mem\[3\]\[124\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_468 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22495_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[45\] _06737_ _06736_ _04945_ _01953_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_90_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24234_ VGND VPWR VPWR VGND clk _00727_ reset_n keymem.key_mem\[11\]\[99\] sky130_fd_sc_hd__dfrtp_2
X_21446_ VGND VPWR VPWR VGND _06184_ _03161_ keymem.key_mem\[5\]\[61\] _06185_ sky130_fd_sc_hd__mux2_2
XFILLER_0_47_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_263_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24165_ VGND VPWR VPWR VGND clk _00658_ reset_n keymem.key_mem\[11\]\[30\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_146_1178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21377_ VGND VPWR _01424_ _06148_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_32_899 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_43_1117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_1128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23116_ VGND VPWR VPWR VGND _07032_ _03479_ keymem.prev_key1_reg\[98\] _07037_ sky130_fd_sc_hd__mux2_2
XFILLER_0_124_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20328_ VGND VPWR VPWR VGND _05580_ _03056_ keymem.key_mem\[9\]\[50\] _05590_ sky130_fd_sc_hd__mux2_2
X_24096_ VGND VPWR VPWR VGND clk _00589_ reset_n keymem.key_mem\[12\]\[89\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_120_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23047_ VGND VPWR VGND VPWR _03789_ key[199] _06995_ _03247_ sky130_fd_sc_hd__a21oi_2
X_20259_ VGND VPWR VPWR VGND _05546_ _11547_ keymem.key_mem\[9\]\[17\] _05554_ sky130_fd_sc_hd__mux2_2
XFILLER_0_228_460 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_21_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14820_ VGND VPWR _00018_ _10285_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_203_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24998_ VGND VPWR VPWR VGND clk _01491_ reset_n keymem.key_mem\[5\]\[95\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_98_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_496 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_235_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_215_187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14751_ VGND VPWR VGND VPWR _10216_ _09665_ _10217_ _09071_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_25_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23949_ VGND VPWR VPWR VGND clk _00442_ reset_n keymem.key_mem\[13\]\[70\] sky130_fd_sc_hd__dfrtp_2
X_11963_ VPWR VGND VGND VPWR _07548_ _07566_ _07532_ sky130_fd_sc_hd__nor2_2
XFILLER_0_98_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_263_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13702_ VGND VPWR _09174_ _09173_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_54_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17470_ VPWR VGND VGND VPWR _03545_ _11021_ _11022_ sky130_fd_sc_hd__nand2_2
X_14682_ VGND VPWR VGND VPWR _08972_ _08999_ _09216_ _09209_ _10149_ sky130_fd_sc_hd__o22a_2
X_11894_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[18\] dec_new_block\[114\]
+ _07511_ sky130_fd_sc_hd__mux2_2
XFILLER_0_131_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_196_573 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16421_ VGND VPWR VPWR VGND _11325_ _11330_ _11222_ _02583_ sky130_fd_sc_hd__or3_2
X_13633_ VGND VPWR _09105_ _09039_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25619_ VGND VPWR VPWR VGND clk _02112_ reset_n keymem.key_mem\[0\]\[76\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_71_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_132_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19140_ VGND VPWR _04928_ _04876_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16352_ VPWR VGND VPWR VGND _02509_ _02514_ _02515_ _02503_ _02506_ sky130_fd_sc_hd__or4b_2
XFILLER_0_183_245 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13564_ VGND VPWR _09036_ _09035_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_27_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_66_284 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_969 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_81_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_211_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15303_ VPWR VGND VGND VPWR _10477_ _10765_ _10440_ sky130_fd_sc_hd__nor2_2
XFILLER_0_26_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12515_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[36\] _07603_ keymem.key_mem\[9\]\[36\]
+ _07592_ _08082_ sky130_fd_sc_hd__a22o_2
X_19071_ VGND VPWR VGND VPWR _04888_ keymem.key_mem_we _10284_ _04878_ _00378_ sky130_fd_sc_hd__a31o_2
X_16283_ VGND VPWR VGND VPWR _11380_ _11253_ _11473_ _11275_ _11412_ _02447_ sky130_fd_sc_hd__o32a_2
X_13495_ VPWR VGND VPWR VGND _08966_ _08948_ _08965_ _08945_ enc_block.block_w2_reg\[1\]
+ _08967_ sky130_fd_sc_hd__a221o_2
XFILLER_0_109_386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_212_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_334 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18022_ VGND VPWR VGND VPWR _03945_ enc_block.round\[3\] _03946_ _00000_ sky130_fd_sc_hd__a21oi_2
X_15234_ VPWR VGND VGND VPWR _10520_ _10697_ _10623_ sky130_fd_sc_hd__nor2_2
X_12446_ VPWR VGND VPWR VGND _08018_ keymem.key_mem\[11\]\[30\] _07809_ keymem.key_mem\[10\]\[30\]
+ _07909_ _08019_ sky130_fd_sc_hd__a221o_2
X_15165_ VGND VPWR _10629_ _10604_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_2_749 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12377_ VPWR VGND VPWR VGND _07955_ keymem.key_mem\[14\]\[24\] _07584_ keymem.key_mem\[6\]\[24\]
+ _07908_ _07956_ sky130_fd_sc_hd__a221o_2
XFILLER_0_22_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_248 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14116_ VPWR VGND VPWR VGND _09587_ _09585_ _09586_ sky130_fd_sc_hd__or2_2
XFILLER_0_142_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15096_ VGND VPWR VGND VPWR _10495_ _10557_ _10488_ _10559_ _10560_ sky130_fd_sc_hd__o22a_2
XFILLER_0_266_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19973_ VPWR VGND VGND VPWR _05402_ _05240_ _05385_ sky130_fd_sc_hd__nand2_2
XFILLER_0_22_398 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18924_ VPWR VGND _04762_ enc_block.block_w0_reg\[9\] enc_block.block_w1_reg\[2\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_14047_ VGND VPWR VPWR VGND _09519_ _08932_ _09517_ _09508_ _09518_ sky130_fd_sc_hd__o31a_2
XFILLER_0_254_717 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_197_1065 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18855_ VPWR VGND VPWR VGND _04700_ _04664_ _04699_ enc_block.block_w2_reg\[10\]
+ _04602_ _00350_ sky130_fd_sc_hd__a221o_2
XFILLER_0_207_655 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17806_ VGND VPWR VGND VPWR _03156_ _03792_ _03795_ _03793_ _03727_ _03800_ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_174_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_98_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18786_ VGND VPWR _04638_ enc_block.block_w3_reg\[20\] enc_block.block_w2_reg\[28\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15998_ VGND VPWR _11453_ _11449_ _11452_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_17737_ VGND VPWR _00176_ _03756_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_253_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14949_ VPWR VGND VPWR VGND _10397_ _10408_ _10403_ _10412_ _10413_ sky130_fd_sc_hd__or4_2
XFILLER_0_210_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17668_ VGND VPWR _00155_ _03708_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19407_ VGND VPWR VGND VPWR _05099_ keymem.key_mem_we _09992_ _05093_ _00503_ sky130_fd_sc_hd__a31o_2
X_16619_ VGND VPWR VPWR VGND _11109_ _02774_ key[28] _02775_ sky130_fd_sc_hd__mux2_2
X_17599_ VGND VPWR VGND VPWR _03657_ _02928_ _02877_ key[126] sky130_fd_sc_hd__o21a_2
XFILLER_0_119_139 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19338_ VGND VPWR VPWR VGND _05046_ _05052_ keymem.key_mem\[13\]\[109\] _05053_ sky130_fd_sc_hd__mux2_2
XFILLER_0_169_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_72_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_2_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_2_Right_170 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19269_ VPWR VGND keymem.key_mem_we _05008_ _03374_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_61_928 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_72_276 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_127_194 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21300_ VGND VPWR _01389_ _06106_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_2_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_356 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22280_ VGND VPWR VPWR VGND _06622_ _03216_ keymem.key_mem\[2\]\[67\] _06629_ sky130_fd_sc_hd__mux2_2
XFILLER_0_72_298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_260_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21231_ VGND VPWR _01356_ _06070_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_79_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_182_1_Right_783 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_142_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21162_ VGND VPWR _01323_ _06034_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20113_ VGND VPWR _00833_ _05475_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_106_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21093_ VGND VPWR _01290_ _05998_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_238_791 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20044_ VGND VPWR _00800_ _05439_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24921_ VGND VPWR VPWR VGND clk _01414_ reset_n keymem.key_mem\[5\]\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_237_290 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_226_975 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_147_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24852_ VGND VPWR VPWR VGND clk _01345_ reset_n keymem.key_mem\[6\]\[77\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_147_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_77_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23803_ VGND VPWR VPWR VGND clk _00296_ reset_n enc_block.block_w0_reg\[22\] sky130_fd_sc_hd__dfrtp_2
X_21995_ VPWR VGND keymem.key_mem\[3\]\[61\] _06478_ _06469_ VPWR VGND sky130_fd_sc_hd__and2_2
X_24783_ VGND VPWR VPWR VGND clk _01276_ reset_n keymem.key_mem\[6\]\[8\] sky130_fd_sc_hd__dfrtp_2
X_20946_ VPWR VGND keymem.key_mem\[7\]\[82\] _05920_ _05899_ VPWR VGND sky130_fd_sc_hd__and2_2
X_23734_ keymem.prev_key0_reg\[90\] clk _00231_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_233_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_152_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_117_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23665_ keymem.prev_key0_reg\[21\] clk _00162_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20877_ VGND VPWR VPWR VGND _05880_ _04955_ keymem.key_mem\[7\]\[50\] _05883_ sky130_fd_sc_hd__mux2_2
XFILLER_0_220_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_230_1368 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25404_ VGND VPWR VPWR VGND clk _01897_ reset_n keymem.key_mem\[2\]\[117\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_796 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22616_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[126\] _06756_ _03793_ _05087_ _02034_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_187_1223 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23596_ VGND VPWR VPWR VGND clk _00097_ reset_n keymem.key_mem\[14\]\[85\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_113_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_906 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_134_1_Left_401 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25335_ VGND VPWR VPWR VGND clk _01828_ reset_n keymem.key_mem\[2\]\[48\] sky130_fd_sc_hd__dfrtp_2
X_22547_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[74\] _06754_ _06753_ _04989_ _01982_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_106_312 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12300_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[18\] _07582_ keymem.key_mem\[8\]\[18\]
+ _07539_ _07885_ sky130_fd_sc_hd__a22o_2
XFILLER_0_49_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13280_ VGND VPWR VGND VPWR _07877_ keymem.key_mem\[10\]\[111\] _08769_ _08771_ _08772_
+ _08020_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_84_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22478_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[33\] _06707_ _06706_ _04922_ _01941_
+ sky130_fd_sc_hd__a22o_2
X_25266_ VGND VPWR VPWR VGND clk _01759_ reset_n keymem.key_mem\[3\]\[107\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_170 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_106_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12231_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[12\] _07645_ _07821_ _07815_ _07822_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_60_961 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21429_ VGND VPWR VPWR VGND _06173_ _03082_ keymem.key_mem\[5\]\[53\] _06176_ sky130_fd_sc_hd__mux2_2
X_24217_ VGND VPWR VPWR VGND clk _00710_ reset_n keymem.key_mem\[11\]\[82\] sky130_fd_sc_hd__dfrtp_2
X_25197_ VGND VPWR VPWR VGND clk _01690_ reset_n keymem.key_mem\[3\]\[38\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_47_1061 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_121_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12162_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[8\] _07578_ keymem.key_mem\[1\]\[8\]
+ _07557_ _07757_ sky130_fd_sc_hd__a22o_2
X_24148_ VGND VPWR VPWR VGND clk _00641_ reset_n keymem.key_mem\[11\]\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_124_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16970_ VPWR VGND VPWR VGND _03098_ _03094_ _03093_ key[183] _03027_ _03099_ sky130_fd_sc_hd__a221o_2
X_12093_ VGND VPWR _07691_ _07690_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24079_ VGND VPWR VPWR VGND clk _00572_ reset_n keymem.key_mem\[12\]\[72\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_21_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15921_ VPWR VGND VGND VPWR _11258_ _11377_ _11286_ sky130_fd_sc_hd__nor2_2
XFILLER_0_21_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_194_1227 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_159_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18640_ VGND VPWR _04507_ enc_block.block_w2_reg\[20\] _04506_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_452 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15852_ VGND VPWR _11308_ _11307_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_614 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_232_934 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_95_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14803_ VGND VPWR VGND VPWR _10267_ _10266_ _10269_ _10268_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_203_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18571_ VGND VPWR _04445_ enc_block.block_w0_reg\[6\] _04444_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15783_ VGND VPWR _11239_ _11238_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12995_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[83\] _07918_ keymem.key_mem\[2\]\[83\]
+ _07697_ _08515_ sky130_fd_sc_hd__a22o_2
XFILLER_0_207_73 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_8_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_1_Left_396 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17522_ VGND VPWR VPWR VGND _09730_ _03589_ key[244] _03590_ sky130_fd_sc_hd__mux2_2
X_14734_ VPWR VGND VGND VPWR _09095_ _10200_ _09136_ sky130_fd_sc_hd__nor2_2
XFILLER_0_52_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_184 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11946_ VPWR VGND VGND VPWR _07548_ _07549_ _07527_ sky130_fd_sc_hd__nor2_2
XFILLER_0_143_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17453_ VGND VPWR VGND VPWR _10828_ _10287_ _03531_ _03530_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_135_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14665_ VGND VPWR VGND VPWR _09333_ _09576_ _09350_ _09423_ _10132_ sky130_fd_sc_hd__o22a_2
X_11877_ VGND VPWR result[105] _07502_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16404_ VPWR VGND VPWR VGND _02563_ _02565_ _02566_ _11578_ _11506_ sky130_fd_sc_hd__or4b_2
XPHY_EDGE_ROW_66_1_Left_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_131_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13616_ VPWR VGND VPWR VGND _09013_ _09004_ _09034_ _08977_ _09088_ sky130_fd_sc_hd__or4_2
X_17384_ VPWR VGND VGND VPWR _03471_ _09630_ _09631_ sky130_fd_sc_hd__nand2_2
X_14596_ VGND VPWR VGND VPWR _09475_ _09423_ _10064_ _09341_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_6_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19123_ VGND VPWR VGND VPWR _04917_ keymem.key_mem_we _02812_ _04908_ _00401_ sky130_fd_sc_hd__a31o_2
XFILLER_0_166_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16335_ VPWR VGND VPWR VGND _02498_ _11255_ _11300_ sky130_fd_sc_hd__or2_2
XFILLER_0_32_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_608 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13547_ VGND VPWR _09019_ _09018_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_67_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_265 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19054_ VGND VPWR _04878_ _04877_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16266_ VPWR VGND VGND VPWR _02417_ _02421_ _02429_ _02430_ sky130_fd_sc_hd__nor3_2
X_13478_ VPWR VGND VPWR VGND _08949_ _08948_ _08946_ _08945_ enc_block.block_w2_reg\[2\]
+ _08950_ sky130_fd_sc_hd__a221o_2
XFILLER_0_67_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_159_2_Left_630 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_259_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18005_ VGND VPWR VGND VPWR _02647_ keymem.prev_key1_reg\[125\] _03679_ _03935_ sky130_fd_sc_hd__a21o_2
X_15217_ VGND VPWR VGND VPWR _10520_ _10510_ _10489_ _10604_ _10680_ sky130_fd_sc_hd__o22a_2
X_12429_ VGND VPWR _08003_ _07744_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16197_ VPWR VGND VPWR VGND _11508_ _11564_ _11290_ _11392_ _02362_ sky130_fd_sc_hd__a22o_2
XFILLER_0_124_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_319 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_471 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_77_12 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15148_ VGND VPWR _10612_ _10611_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_22_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_579 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_26_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_267_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_142_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1138 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15079_ VGND VPWR _10543_ _10441_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_103_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19956_ VGND VPWR VPWR VGND _05389_ _09992_ keymem.key_mem\[10\]\[3\] _05393_ sky130_fd_sc_hd__mux2_2
XFILLER_0_177_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18907_ VPWR VGND VGND VPWR _04747_ _04684_ _04746_ sky130_fd_sc_hd__nand2_2
XFILLER_0_103_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19887_ VGND VPWR VPWR VGND _05350_ keymem.key_mem\[11\]\[100\] _03492_ _05355_ sky130_fd_sc_hd__mux2_2
XFILLER_0_177_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18838_ VGND VPWR _04685_ _04606_ _04684_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_945 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_179_315 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_117_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18769_ VPWR VGND VGND VPWR _04613_ _04623_ _04005_ sky130_fd_sc_hd__nor2_2
XFILLER_0_250_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_179_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_218_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20800_ VGND VPWR VGND VPWR _05841_ keymem.key_mem_we _11099_ _05838_ _01154_ sky130_fd_sc_hd__a31o_2
X_21780_ VGND VPWR VPWR VGND _06355_ _03426_ keymem.key_mem\[4\]\[91\] _06361_ sky130_fd_sc_hd__mux2_2
XFILLER_0_114_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20731_ VGND VPWR VPWR VGND _05794_ _03573_ keymem.key_mem\[8\]\[113\] _05802_ sky130_fd_sc_hd__mux2_2
XFILLER_0_153_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23450_ VPWR VGND _07316_ _07315_ enc_block.round_key\[25\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_114_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20662_ VGND VPWR VPWR VGND _05761_ _03329_ keymem.key_mem\[8\]\[80\] _05766_ sky130_fd_sc_hd__mux2_2
XFILLER_0_188_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_133_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22401_ VGND VPWR VPWR VGND _06553_ _03654_ keymem.key_mem\[2\]\[125\] _06692_ sky130_fd_sc_hd__mux2_2
XFILLER_0_162_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23381_ VPWR VGND VGND VPWR _07192_ _07255_ _04169_ sky130_fd_sc_hd__nor2_2
X_20593_ VGND VPWR VPWR VGND _05725_ _03024_ keymem.key_mem\[8\]\[47\] _05730_ sky130_fd_sc_hd__mux2_2
XFILLER_0_2_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_2_Right_171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25120_ VGND VPWR VPWR VGND clk _01613_ reset_n keymem.key_mem\[4\]\[89\] sky130_fd_sc_hd__dfrtp_2
X_22332_ VGND VPWR VPWR VGND _06647_ _03434_ keymem.key_mem\[2\]\[92\] _06656_ sky130_fd_sc_hd__mux2_2
XFILLER_0_264_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_950 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25051_ VGND VPWR VPWR VGND clk _01544_ reset_n keymem.key_mem\[4\]\[20\] sky130_fd_sc_hd__dfrtp_2
X_22263_ VGND VPWR VPWR VGND _06611_ _03139_ keymem.key_mem\[2\]\[59\] _06620_ sky130_fd_sc_hd__mux2_2
XFILLER_0_103_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24002_ VGND VPWR VPWR VGND clk _00495_ reset_n keymem.key_mem\[13\]\[123\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_44_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21214_ VGND VPWR _01348_ _06061_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22194_ VGND VPWR VPWR VGND _06578_ _02742_ keymem.key_mem\[2\]\[26\] _06584_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_183_1_Right_784 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_125_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_2_Left_551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21145_ VGND VPWR _01315_ _06025_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_111_381 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_22_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_10_891 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_121_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21076_ VGND VPWR _01282_ _05989_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_22_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20027_ VGND VPWR _00792_ _05430_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24904_ VGND VPWR VPWR VGND clk _01397_ reset_n keymem.key_mem\[5\]\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_236_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24835_ VGND VPWR VPWR VGND clk _01328_ reset_n keymem.key_mem\[6\]\[60\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_236_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_240_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11800_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[3\] dec_new_block\[67\]
+ _07464_ sky130_fd_sc_hd__mux2_2
X_12780_ VGND VPWR VGND VPWR _08322_ _07753_ keymem.key_mem\[8\]\[61\] _08319_ _08321_
+ sky130_fd_sc_hd__a211o_2
X_24766_ VGND VPWR VPWR VGND clk _01259_ reset_n keymem.key_mem\[7\]\[119\] sky130_fd_sc_hd__dfrtp_2
X_21978_ VGND VPWR VGND VPWR _06468_ keymem.key_mem_we _03083_ _06446_ _01705_ sky130_fd_sc_hd__a31o_2
X_11731_ VGND VPWR result[32] _07429_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_132_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23717_ keymem.prev_key0_reg\[73\] clk _00214_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20929_ VGND VPWR _01214_ _05910_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24697_ VGND VPWR VPWR VGND clk _01190_ reset_n keymem.key_mem\[7\]\[50\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_260_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14450_ VGND VPWR _09918_ _09336_ _09919_ _09396_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_49_582 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_132_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_22_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11662_ VGND VPWR VGND VPWR _00008_ _07393_ enc_block.enc_ctrl_reg\[3\] _07395_ enc_block.enc_ctrl_reg\[2\]
+ sky130_fd_sc_hd__a211o_2
X_23648_ keymem.prev_key0_reg\[4\] clk _00145_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_13401_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[123\] _07560_ keymem.key_mem\[1\]\[123\]
+ _07556_ _08881_ sky130_fd_sc_hd__a22o_2
XFILLER_0_14_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14381_ VGND VPWR VGND VPWR _09850_ _09827_ _09240_ _09851_ sky130_fd_sc_hd__a21o_2
XFILLER_0_52_714 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23579_ VGND VPWR VPWR VGND clk _00080_ reset_n keymem.key_mem\[14\]\[68\] sky130_fd_sc_hd__dfrtp_2
X_16120_ VGND VPWR _11573_ _11211_ _11574_ _11420_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_64_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_153_259 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_88_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25318_ VGND VPWR VPWR VGND clk _01811_ reset_n keymem.key_mem\[2\]\[31\] sky130_fd_sc_hd__dfrtp_2
X_13332_ VPWR VGND VPWR VGND _08818_ keymem.key_mem\[3\]\[116\] _07690_ keymem.key_mem\[12\]\[116\]
+ _07788_ _08819_ sky130_fd_sc_hd__a221o_2
XFILLER_0_91_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16051_ VPWR VGND VGND VPWR _11469_ _11506_ _11367_ sky130_fd_sc_hd__nor2_2
XFILLER_0_45_1009 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_243_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25249_ VGND VPWR VPWR VGND clk _01742_ reset_n keymem.key_mem\[3\]\[90\] sky130_fd_sc_hd__dfrtp_2
X_13263_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[109\] _07621_ keymem.key_mem\[8\]\[109\]
+ _07929_ _08757_ sky130_fd_sc_hd__a22o_2
XFILLER_0_161_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_106_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_460 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15002_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[11\] _08989_ _10466_ _08983_ _10406_
+ _10407_ sky130_fd_sc_hd__a32oi_2
X_12214_ VGND VPWR enc_block.round_key\[11\] _07805_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13194_ VGND VPWR VGND VPWR _07793_ keymem.key_mem\[0\]\[102\] _08694_ _08689_ _08687_
+ _08695_ sky130_fd_sc_hd__o32a_2
XFILLER_0_121_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_666 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19810_ VGND VPWR VPWR VGND _05314_ keymem.key_mem\[11\]\[63\] _03184_ _05315_ sky130_fd_sc_hd__mux2_2
X_12145_ VPWR VGND VPWR VGND _07740_ keymem.key_mem\[6\]\[7\] _07739_ keymem.key_mem\[9\]\[7\]
+ _07738_ _07741_ sky130_fd_sc_hd__a221o_2
XFILLER_0_47_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_739 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16953_ VGND VPWR _03084_ _09863_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19741_ VGND VPWR _00658_ _05278_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12076_ VPWR VGND VPWR VGND _07675_ keymem.key_mem\[9\]\[3\] _07672_ keymem.key_mem\[1\]\[3\]
+ _07671_ _07676_ sky130_fd_sc_hd__a221o_2
X_15904_ VPWR VGND VPWR VGND _11265_ _11248_ _11243_ _11166_ _11360_ sky130_fd_sc_hd__or4_2
X_19672_ VGND VPWR VPWR VGND keymem.round_ctr_reg\[2\] _05240_ keymem.round_ctr_reg\[3\]
+ sky130_fd_sc_hd__and2b_2
X_16884_ VGND VPWR VGND VPWR _03021_ _09721_ _09795_ key[47] sky130_fd_sc_hd__o21a_2
X_18623_ VPWR VGND VGND VPWR _04491_ _04492_ _04478_ sky130_fd_sc_hd__nor2_2
XFILLER_0_159_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15835_ VPWR VGND VGND VPWR _11266_ _11291_ _11167_ sky130_fd_sc_hd__nor2_2
XFILLER_0_204_433 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_232_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_231_241 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18554_ VPWR VGND VGND VPWR _04429_ _04430_ _04077_ sky130_fd_sc_hd__nor2_2
X_15766_ VGND VPWR _11222_ _11221_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_59_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_937 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12978_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[81\] _08090_ keymem.key_mem\[2\]\[81\]
+ _08131_ _08500_ sky130_fd_sc_hd__a22o_2
X_17505_ VGND VPWR VPWR VGND _10366_ _11622_ key[114] _03575_ sky130_fd_sc_hd__mux2_2
X_14717_ VPWR VGND VGND VPWR _09075_ _10182_ _10183_ _10184_ sky130_fd_sc_hd__nor3_2
X_18485_ _04366_ _04368_ _04294_ _04367_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_11929_ VPWR VGND VGND VPWR _07532_ _07525_ _07526_ sky130_fd_sc_hd__nand2_2
X_15697_ _10552_ _11153_ keymem.prev_key1_reg\[112\] _10652_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_200_650 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17436_ VGND VPWR VGND VPWR _03516_ _03515_ _03514_ _10092_ sky130_fd_sc_hd__o21a_2
XFILLER_0_137_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14648_ VPWR VGND VGND VPWR _09559_ _09368_ _09343_ _10115_ sky130_fd_sc_hd__nor3_2
XFILLER_0_200_683 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17367_ VGND VPWR VGND VPWR key[95] _09930_ _03455_ _03454_ _03456_ sky130_fd_sc_hd__o22a_2
X_14579_ VPWR VGND VGND VPWR _09383_ _10047_ _09576_ sky130_fd_sc_hd__nor2_2
XFILLER_0_3_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19106_ VGND VPWR _04908_ _04877_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_6_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_67_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16318_ VGND VPWR _00032_ _02481_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_103_86 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_15_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17298_ VGND VPWR _00099_ _03394_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19037_ VGND VPWR _04863_ _04657_ _04862_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16249_ VPWR VGND VPWR VGND _11508_ _11564_ _11290_ _11503_ _02413_ sky130_fd_sc_hd__a22o_2
XFILLER_0_203_1009 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_514 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_396 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_227_547 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_255_867 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19939_ VGND VPWR VPWR VGND _05372_ keymem.key_mem\[11\]\[125\] _03654_ _05382_ sky130_fd_sc_hd__mux2_2
XFILLER_0_177_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22950_ VGND VPWR _02208_ _06937_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_78_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21901_ VGND VPWR _06427_ _06405_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_74_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22881_ VGND VPWR VGND VPWR _02182_ _06894_ _06882_ keymem.prev_key1_reg\[5\] sky130_fd_sc_hd__o21a_2
XFILLER_0_39_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24620_ VGND VPWR VPWR VGND clk _01113_ reset_n keymem.key_mem\[8\]\[101\] sky130_fd_sc_hd__dfrtp_2
X_21832_ VGND VPWR _06388_ _06258_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_37_1060 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_214_1149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_190_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21763_ VGND VPWR VPWR VGND _06344_ _03355_ keymem.key_mem\[4\]\[83\] _06352_ sky130_fd_sc_hd__mux2_2
X_24551_ VGND VPWR VPWR VGND clk _01044_ reset_n keymem.key_mem\[8\]\[32\] sky130_fd_sc_hd__dfrtp_2
X_23502_ VPWR VGND VGND VPWR _07361_ _07362_ enc_block.round_key\[31\] sky130_fd_sc_hd__nor2_2
X_20714_ VGND VPWR VPWR VGND _05783_ _03525_ keymem.key_mem\[8\]\[105\] _05793_ sky130_fd_sc_hd__mux2_2
X_24482_ VGND VPWR VPWR VGND clk _00975_ reset_n keymem.key_mem\[9\]\[91\] sky130_fd_sc_hd__dfrtp_2
X_21694_ VGND VPWR VPWR VGND _06308_ _03056_ keymem.key_mem\[4\]\[50\] _06316_ sky130_fd_sc_hd__mux2_2
XFILLER_0_65_349 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_114_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_384 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23433_ VGND VPWR VGND VPWR _07299_ _07298_ _07301_ _07297_ sky130_fd_sc_hd__a21oi_2
X_20645_ VGND VPWR VPWR VGND _05747_ _03259_ keymem.key_mem\[8\]\[72\] _05757_ sky130_fd_sc_hd__mux2_2
XFILLER_0_11_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_179 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_230_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23364_ VPWR VGND _07239_ _07176_ _07166_ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_85_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20576_ VGND VPWR VPWR VGND _05714_ _02945_ keymem.key_mem\[8\]\[39\] _05721_ sky130_fd_sc_hd__mux2_2
XFILLER_0_149_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25103_ VGND VPWR VPWR VGND clk _01596_ reset_n keymem.key_mem\[4\]\[72\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_85_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22315_ VGND VPWR _06647_ _06552_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23295_ VGND VPWR _07177_ _07099_ _07176_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_791 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22246_ VGND VPWR _06611_ _06553_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25034_ VGND VPWR VPWR VGND clk _01527_ reset_n keymem.key_mem\[4\]\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_239_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22177_ VGND VPWR VPWR VGND _06565_ _02339_ keymem.key_mem\[2\]\[18\] _06575_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_184_1_Right_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21128_ VGND VPWR _01307_ _06016_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_258_1032 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_255_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_219_1016 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13950_ VGND VPWR _09422_ _09421_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_233_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21059_ VGND VPWR VPWR VGND _05972_ _10369_ keymem.key_mem\[6\]\[7\] _05980_ sky130_fd_sc_hd__mux2_2
XFILLER_0_96_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12901_ VGND VPWR enc_block.round_key\[73\] _08430_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13881_ VGND VPWR _09353_ _09352_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_9_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15620_ VGND VPWR VGND VPWR _10618_ _10546_ _10441_ _11078_ sky130_fd_sc_hd__a21o_2
XFILLER_0_57_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24818_ VGND VPWR VPWR VGND clk _01311_ reset_n keymem.key_mem\[6\]\[43\] sky130_fd_sc_hd__dfrtp_2
X_12832_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[67\] _07759_ keymem.key_mem\[11\]\[67\]
+ _07761_ _08368_ sky130_fd_sc_hd__a22o_2
XFILLER_0_9_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_110 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25798_ keymem.prev_key1_reg\[114\] clk _02291_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_202_959 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_806 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15551_ VGND VPWR VGND VPWR _11009_ _11007_ _11010_ _10705_ _10549_ sky130_fd_sc_hd__nand4_2
XFILLER_0_9_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12763_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[60\] _07695_ keymem.key_mem\[14\]\[60\]
+ _08003_ _08306_ sky130_fd_sc_hd__a22o_2
X_24749_ VGND VPWR VPWR VGND clk _01242_ reset_n keymem.key_mem\[7\]\[102\] sky130_fd_sc_hd__dfrtp_2
X_14502_ VGND VPWR VGND VPWR _09969_ _09181_ _09971_ _09970_ sky130_fd_sc_hd__a21oi_2
X_18270_ VPWR VGND VGND VPWR _04174_ _04089_ _04173_ sky130_fd_sc_hd__nand2_2
X_11714_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[24\] dec_new_block\[24\]
+ _07421_ sky130_fd_sc_hd__mux2_2
X_15482_ VGND VPWR VGND VPWR _10574_ _10482_ _10508_ _10942_ sky130_fd_sc_hd__a21o_2
X_12694_ VGND VPWR VGND VPWR _07808_ keymem.key_mem\[12\]\[53\] _08240_ _08242_ _08244_
+ _08243_ sky130_fd_sc_hd__a2111o_2
XPHY_EDGE_ROW_253_Right_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17221_ VGND VPWR VGND VPWR _11441_ keymem.prev_key0_reg\[80\] _03325_ _10327_ sky130_fd_sc_hd__nand3_2
X_14433_ VPWR VGND VGND VPWR _09902_ _09900_ _09901_ sky130_fd_sc_hd__nand2_2
X_11645_ VPWR VGND VGND VPWR _07383_ init keymem.key_mem_ctrl_reg\[0\] sky130_fd_sc_hd__nand2_2
XFILLER_0_140_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_167_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17152_ VPWR VGND VPWR VGND _03263_ keymem.prev_key0_reg\[73\] sky130_fd_sc_hd__inv_2
X_14364_ VPWR VGND VGND VPWR _09834_ _09832_ _09833_ sky130_fd_sc_hd__nand2_2
XFILLER_0_52_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_68_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_167_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_909 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_91_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16103_ VGND VPWR VGND VPWR _09511_ _11555_ _11553_ _11554_ _11557_ sky130_fd_sc_hd__a31o_2
XFILLER_0_247_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13315_ VGND VPWR enc_block.round_key\[114\] _08803_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17083_ VPWR VGND VPWR VGND _03201_ _03199_ _03198_ key[193] _03027_ _03202_ sky130_fd_sc_hd__a221o_2
X_14295_ VPWR VGND VGND VPWR _09441_ _09765_ _09380_ sky130_fd_sc_hd__nor2_2
XFILLER_0_29_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16034_ VGND VPWR VPWR VGND _11487_ _11488_ _11486_ _11489_ sky130_fd_sc_hd__or3_2
X_13246_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[107\] _08714_ _08741_ _08737_ _08742_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_0_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13177_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[101\] _07685_ keymem.key_mem\[1\]\[101\]
+ _07624_ _08679_ sky130_fd_sc_hd__a22o_2
XFILLER_0_249_694 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_631 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_229_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12128_ VGND VPWR _07725_ _07724_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17985_ VGND VPWR VPWR VGND _03674_ _03921_ keymem.prev_key0_reg\[118\] _03922_ sky130_fd_sc_hd__mux2_2
XFILLER_0_178_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1086 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_139_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16936_ VGND VPWR VPWR VGND _02986_ keymem.key_mem\[14\]\[51\] _03068_ _03069_ sky130_fd_sc_hd__mux2_2
XFILLER_0_263_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12059_ VGND VPWR _07659_ _07595_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19724_ VGND VPWR _00650_ _05269_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_178_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_75_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16867_ VPWR VGND VPWR VGND _03005_ _03001_ _03000_ key[173] _02875_ _03006_ sky130_fd_sc_hd__a221o_2
XFILLER_0_254_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19655_ VGND VPWR _00619_ _05231_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_219_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_75_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15818_ VGND VPWR VPWR VGND _11272_ _11273_ _11226_ _11274_ sky130_fd_sc_hd__or3_2
X_18606_ VPWR VGND VGND VPWR _04380_ _04477_ _04169_ sky130_fd_sc_hd__nor2_2
XFILLER_0_254_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19586_ VGND VPWR _00586_ _05195_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16798_ VPWR VGND VGND VPWR _02943_ _11456_ _10317_ sky130_fd_sc_hd__nand2_2
X_18537_ VPWR VGND VGND VPWR _04380_ _04415_ _04095_ sky130_fd_sc_hd__nor2_2
XFILLER_0_215_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15749_ VGND VPWR _11205_ _11204_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_133_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_914 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18468_ VGND VPWR _04352_ enc_block.block_w1_reg\[27\] enc_block.block_w1_reg\[31\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_7_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17419_ VPWR VGND VGND VPWR _03501_ _10263_ _10264_ sky130_fd_sc_hd__nand2_2
X_18399_ VGND VPWR _04291_ _03950_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_184_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_12_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_371 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_522 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20430_ VGND VPWR _00982_ _05643_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_172_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_146_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_125_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20361_ VGND VPWR _00949_ _05607_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_226_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22100_ VGND VPWR VPWR VGND _06527_ _05056_ keymem.key_mem\[3\]\[111\] _06533_ sky130_fd_sc_hd__mux2_2
X_23080_ VGND VPWR _02260_ _07015_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_222_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20292_ VGND VPWR _00916_ _05571_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_2_162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22031_ VGND VPWR VPWR VGND _06494_ _04997_ keymem.key_mem\[3\]\[78\] _06497_ sky130_fd_sc_hd__mux2_2
XFILLER_0_41_1215 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_80_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_496 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_100_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_122_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23982_ VGND VPWR VPWR VGND clk _00475_ reset_n keymem.key_mem\[13\]\[103\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_143_1_Left_410 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25721_ keymem.prev_key1_reg\[37\] clk _02214_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_78_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22933_ VPWR VGND VPWR VGND _06927_ keymem.prev_key1_reg\[25\] _06926_ sky130_fd_sc_hd__or2_2
XFILLER_0_155_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1166 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_233_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25652_ VGND VPWR VPWR VGND clk _02145_ reset_n keymem.key_mem\[0\]\[109\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22864_ VGND VPWR _06882_ _06881_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_64_90 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24603_ VGND VPWR VPWR VGND clk _01096_ reset_n keymem.key_mem\[8\]\[84\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_233_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21815_ VGND VPWR _01631_ _06379_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_6_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25583_ VGND VPWR VPWR VGND clk _02076_ reset_n keymem.key_mem\[0\]\[40\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_151_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22795_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[98\] _06850_ _06849_ _05029_ _02134_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_65_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24534_ VGND VPWR VPWR VGND clk _01027_ reset_n keymem.key_mem\[8\]\[15\] sky130_fd_sc_hd__dfrtp_2
X_21746_ VPWR VGND VGND VPWR _06259_ _06343_ keymem.key_mem\[4\]\[75\] sky130_fd_sc_hd__nor2_2
XFILLER_0_241_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24465_ VGND VPWR VPWR VGND clk _00958_ reset_n keymem.key_mem\[9\]\[74\] sky130_fd_sc_hd__dfrtp_2
X_21677_ VGND VPWR VPWR VGND _06297_ _02972_ keymem.key_mem\[4\]\[42\] _06307_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_382 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23416_ VPWR VGND VPWR VGND _07286_ _07211_ _07284_ sky130_fd_sc_hd__or2_2
XFILLER_0_34_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20628_ VGND VPWR _01075_ _05748_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24396_ VGND VPWR VPWR VGND clk _00889_ reset_n keymem.key_mem\[9\]\[5\] sky130_fd_sc_hd__dfrtp_2
X_23347_ VPWR VGND VGND VPWR _07224_ _07148_ _07223_ sky130_fd_sc_hd__nand2_2
X_20559_ VGND VPWR VPWR VGND _05703_ _02861_ keymem.key_mem\[8\]\[31\] _05712_ sky130_fd_sc_hd__mux2_2
X_13100_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[93\] _07984_ keymem.key_mem\[4\]\[93\]
+ _08077_ _08610_ sky130_fd_sc_hd__a22o_2
X_14080_ _09550_ _09551_ _09463_ _09364_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_23278_ _07160_ _07162_ _04103_ _07161_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_14_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13031_ VGND VPWR VGND VPWR _08548_ _07580_ keymem.key_mem\[12\]\[86\] _08545_ _08547_
+ sky130_fd_sc_hd__a211o_2
X_25017_ VGND VPWR VPWR VGND clk _01510_ reset_n keymem.key_mem\[5\]\[114\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_162_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22229_ VGND VPWR _01822_ _06602_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_106_2_Left_577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_119_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_185_1_Right_786 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_218_355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_75_1_Left_342 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_219_889 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17770_ VGND VPWR VPWR VGND _03763_ _03043_ keymem.prev_key0_reg\[49\] _03776_ sky130_fd_sc_hd__mux2_2
XFILLER_0_234_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14982_ VPWR VGND VPWR VGND _10424_ _10445_ _10444_ _10443_ _10446_ sky130_fd_sc_hd__or4_2
X_16721_ VGND VPWR VGND VPWR _02873_ _02868_ _02865_ _02871_ _02872_ sky130_fd_sc_hd__a211o_2
X_13933_ VGND VPWR VGND VPWR _09399_ _09349_ _09404_ _09401_ _09405_ sky130_fd_sc_hd__o22a_2
XFILLER_0_57_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19440_ VGND VPWR VGND VPWR _05117_ keymem.key_mem_we _02340_ _05109_ _00518_ sky130_fd_sc_hd__a31o_2
X_16652_ _02804_ _02807_ _02803_ _02805_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_18_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13864_ VGND VPWR _09336_ _09335_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_92_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15603_ VGND VPWR VGND VPWR _10635_ _10441_ _11061_ _10476_ sky130_fd_sc_hd__a21oi_2
X_12815_ VGND VPWR VGND VPWR _07542_ keymem.key_mem\[8\]\[65\] _08350_ _08352_ _08353_
+ _08243_ sky130_fd_sc_hd__a2111o_2
X_19371_ VPWR VGND keymem.key_mem_we _05075_ _03620_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_215_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16583_ VPWR VGND VPWR VGND _02741_ _10325_ _02738_ _02739_ _02740_ _10281_ sky130_fd_sc_hd__o311a_2
X_13795_ VGND VPWR VPWR VGND _09261_ _09266_ _09254_ _09267_ sky130_fd_sc_hd__or3_2
XFILLER_0_202_778 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_316 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18322_ VPWR VGND _04222_ _04221_ enc_block.round_key\[118\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_210_1300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15534_ VPWR VGND VPWR VGND _10983_ _10992_ _10987_ _10493_ _10993_ sky130_fd_sc_hd__or4_2
XFILLER_0_56_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_210_1311 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12746_ VGND VPWR VGND VPWR _07842_ keymem.key_mem\[9\]\[58\] _08288_ _08290_ _08291_
+ _08020_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_60_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18253_ VPWR VGND VPWR VGND _04159_ _03970_ _11439_ sky130_fd_sc_hd__or2_2
XFILLER_0_70_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15465_ VPWR VGND VGND VPWR _10566_ _10925_ _10569_ sky130_fd_sc_hd__nor2_2
X_12677_ VGND VPWR VGND VPWR _08229_ _08150_ keymem.key_mem\[3\]\[51\] _08226_ _08228_
+ sky130_fd_sc_hd__a211o_2
X_17204_ VGND VPWR VPWR VGND _02864_ _11092_ keymem.prev_key0_reg\[78\] _03310_ sky130_fd_sc_hd__or3_2
X_14416_ VGND VPWR VGND VPWR _09780_ _09364_ _09776_ _09884_ _09885_ _09602_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_25_522 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_61 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18184_ VPWR VGND VGND VPWR _04095_ _04096_ _04041_ sky130_fd_sc_hd__nor2_2
XFILLER_0_154_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11628_ VGND VPWR VGND VPWR aes_core_ctrl_reg\[2\] keymem.ready _07369_ _07368_ sky130_fd_sc_hd__a21oi_2
X_15396_ VGND VPWR VGND VPWR _10538_ _10668_ _10489_ _10547_ _10857_ sky130_fd_sc_hd__o22a_2
XFILLER_0_52_341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_68_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17135_ VGND VPWR VGND VPWR _03248_ keymem.prev_key0_reg\[71\] _10364_ _10363_ _09988_
+ sky130_fd_sc_hd__o211ai_2
X_14347_ VGND VPWR VGND VPWR _09107_ _09174_ _09134_ _09149_ _09817_ sky130_fd_sc_hd__o22a_2
XFILLER_0_68_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17066_ VGND VPWR _00075_ _03186_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_180_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14278_ VGND VPWR VGND VPWR _09392_ _09389_ _09456_ _09404_ _09748_ sky130_fd_sc_hd__o22a_2
XFILLER_0_257_918 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_229_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_208_1295 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16017_ VPWR VGND VGND VPWR _11472_ _11470_ _11471_ sky130_fd_sc_hd__nand2_2
X_13229_ VPWR VGND VPWR VGND _08725_ keymem.key_mem\[6\]\[106\] _07739_ keymem.key_mem\[4\]\[106\]
+ _07637_ _08726_ sky130_fd_sc_hd__a221o_2
XFILLER_0_180_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1440 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17968_ VGND VPWR VPWR VGND _03876_ key[241] keymem.prev_key1_reg\[113\] _03910_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_85_89 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_139_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_100_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19707_ VGND VPWR VPWR VGND _05259_ keymem.key_mem\[11\]\[14\] _11099_ _05261_ sky130_fd_sc_hd__mux2_2
X_16919_ VPWR VGND VPWR VGND keymem.prev_key1_reg\[50\] _03053_ _11556_ _11557_ sky130_fd_sc_hd__or3b_2
XFILLER_0_224_358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_79_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17899_ VGND VPWR VGND VPWR _03863_ keymem.prev_key0_reg\[90\] _00231_ _03736_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_174_1269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_36_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19638_ VGND VPWR _00611_ _05222_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_192_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_215_1255 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19569_ VGND VPWR _00578_ _05186_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_149_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21600_ VGND VPWR VPWR VGND _06263_ _10193_ keymem.key_mem\[4\]\[5\] _06267_ sky130_fd_sc_hd__mux2_2
X_22580_ VGND VPWR VPWR VGND _06701_ keymem.key_mem\[1\]\[95\] _03460_ _06773_ sky130_fd_sc_hd__mux2_2
XFILLER_0_220_597 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_850 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_145_310 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21531_ VGND VPWR VPWR VGND _06220_ _03506_ keymem.key_mem\[5\]\[102\] _06229_ sky130_fd_sc_hd__mux2_2
XFILLER_0_157_192 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21462_ VGND VPWR VPWR VGND _06184_ _03234_ keymem.key_mem\[5\]\[69\] _06193_ sky130_fd_sc_hd__mux2_2
X_24250_ VGND VPWR VPWR VGND clk _00743_ reset_n keymem.key_mem\[11\]\[115\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_141_72 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_86_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23201_ VGND VPWR VGND VPWR _00001_ _07381_ _07092_ _03949_ sky130_fd_sc_hd__a21oi_2
X_20413_ VGND VPWR _00974_ _05634_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24181_ VGND VPWR VPWR VGND clk _00674_ reset_n keymem.key_mem\[11\]\[46\] sky130_fd_sc_hd__dfrtp_2
X_21393_ VGND VPWR VPWR VGND _06151_ _02913_ keymem.key_mem\[5\]\[36\] _06157_ sky130_fd_sc_hd__mux2_2
XFILLER_0_47_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23132_ VGND VPWR VPWR VGND _07032_ _07046_ keymem.prev_key1_reg\[104\] _07047_ sky130_fd_sc_hd__mux2_2
X_20344_ VGND VPWR _00941_ _05598_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23063_ VGND VPWR VGND VPWR _07005_ _03303_ _03301_ _03305_ _06951_ sky130_fd_sc_hd__a211o_2
XFILLER_0_109_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20275_ VGND VPWR _00908_ _05562_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22014_ VGND VPWR VPWR VGND _06462_ _04983_ keymem.key_mem\[3\]\[70\] _06488_ sky130_fd_sc_hd__mux2_2
XFILLER_0_243_601 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_243_623 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_157_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23965_ VGND VPWR VPWR VGND clk _00458_ reset_n keymem.key_mem\[13\]\[86\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25704_ keymem.prev_key1_reg\[20\] clk _02197_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22916_ VGND VPWR _02196_ _06915_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_19_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23896_ VGND VPWR VPWR VGND clk _00389_ reset_n keymem.key_mem\[13\]\[17\] sky130_fd_sc_hd__dfrtp_2
X_25635_ VGND VPWR VPWR VGND clk _02128_ reset_n keymem.key_mem\[0\]\[92\] sky130_fd_sc_hd__dfrtp_2
X_22847_ VPWR VGND VPWR VGND _06871_ keymem.key_mem_we keymem.round_ctr_reg\[0\] sky130_fd_sc_hd__or2_2
X_12600_ VPWR VGND VPWR VGND _08158_ keymem.key_mem\[5\]\[44\] _07683_ keymem.key_mem\[4\]\[44\]
+ _07637_ _08159_ sky130_fd_sc_hd__a221o_2
X_13580_ VGND VPWR VPWR VGND _09010_ _09051_ _09009_ _09052_ sky130_fd_sc_hd__or3_2
X_25566_ VGND VPWR VPWR VGND clk _02059_ reset_n keymem.key_mem\[0\]\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22778_ VGND VPWR VPWR VGND _06784_ keymem.key_mem\[0\]\[87\] _03393_ _06851_ sky130_fd_sc_hd__mux2_2
XFILLER_0_136_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24517_ VGND VPWR VPWR VGND clk _01010_ reset_n keymem.key_mem\[9\]\[126\] sky130_fd_sc_hd__dfrtp_2
X_12531_ VGND VPWR _08096_ _08052_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21729_ VGND VPWR _01590_ _06334_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_53_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25497_ VGND VPWR VPWR VGND clk _01990_ reset_n keymem.key_mem\[1\]\[82\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_87_1226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15250_ VPWR VGND VPWR VGND _10704_ _10712_ _10707_ _10700_ _10713_ sky130_fd_sc_hd__or4_2
XFILLER_0_129_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_19_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24448_ VGND VPWR VPWR VGND clk _00941_ reset_n keymem.key_mem\[9\]\[57\] sky130_fd_sc_hd__dfrtp_2
X_12462_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[31\] _07639_ keymem.key_mem\[11\]\[31\]
+ _07599_ _08034_ sky130_fd_sc_hd__a22o_2
XFILLER_0_168_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14201_ VPWR VGND VGND VPWR _09134_ _09672_ _09080_ sky130_fd_sc_hd__nor2_2
XFILLER_0_129_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15181_ VPWR VGND VPWR VGND _10457_ _10644_ _10430_ _10419_ _10645_ sky130_fd_sc_hd__or4_2
XFILLER_0_35_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12393_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[25\] _07568_ keymem.key_mem\[2\]\[25\]
+ _07732_ _07971_ sky130_fd_sc_hd__a22o_2
X_24379_ VGND VPWR VPWR VGND clk _00872_ reset_n keymem.key_mem\[10\]\[116\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_22_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14132_ _09363_ _09603_ _09550_ _09553_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_266_704 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_238_406 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_205_1446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_39_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18940_ VPWR VGND _04777_ _04776_ enc_block.round_key\[51\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_14063_ VGND VPWR VGND VPWR _09535_ _09519_ _09514_ _09534_ _09532_ _09509_ sky130_fd_sc_hd__a32o_2
XFILLER_0_162_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_123_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13014_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[85\] _07743_ keymem.key_mem\[8\]\[85\]
+ _07958_ _08532_ sky130_fd_sc_hd__a22o_2
X_18871_ VPWR VGND VPWR VGND _04714_ block[44] _04576_ enc_block.block_w0_reg\[12\]
+ _04666_ _04715_ sky130_fd_sc_hd__a221o_2
XFILLER_0_218_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_206_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17822_ VGND VPWR VPWR VGND _03719_ key[195] keymem.prev_key1_reg\[67\] _03810_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_186_1_Right_787 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_55_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14965_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[14\] _08955_ _10429_ _08942_ _10427_
+ _10428_ sky130_fd_sc_hd__a32oi_2
X_17753_ VGND VPWR VPWR VGND _03719_ key[170] keymem.prev_key1_reg\[42\] _03766_ sky130_fd_sc_hd__mux2_2
XFILLER_0_136_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_998 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_226_50 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13916_ VGND VPWR _09388_ _09387_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16704_ _02855_ _02857_ _02854_ _02856_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_17684_ VGND VPWR _03719_ _03211_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_226_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14896_ VGND VPWR VGND VPWR _10359_ _10336_ _10360_ _10361_ sky130_fd_sc_hd__a21o_2
XFILLER_0_216_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_210 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19423_ VGND VPWR VPWR VGND _05092_ _04894_ keymem.key_mem\[12\]\[11\] _05108_ sky130_fd_sc_hd__mux2_2
X_16635_ VGND VPWR VGND VPWR _02536_ keymem.rcon_logic.tmp_rcon\[6\] _02790_ _11301_
+ sky130_fd_sc_hd__nand3_2
X_13847_ VGND VPWR _09319_ _09254_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_202_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_29_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_69_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19354_ VGND VPWR _00486_ _05063_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16566_ VGND VPWR VGND VPWR _11618_ _11589_ keymem.rcon_reg\[2\] _02724_ sky130_fd_sc_hd__a21o_2
X_13778_ enc_block.sword_ctr_reg\[1\] _09250_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[27\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_71_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18305_ _04204_ _04206_ _04203_ _04205_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_15517_ VGND VPWR _10977_ _10976_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19285_ VPWR VGND keymem.key_mem\[13\]\[91\] _05018_ _04879_ VPWR VGND sky130_fd_sc_hd__and2_2
X_12729_ VPWR VGND VPWR VGND _08275_ keymem.key_mem\[5\]\[56\] _08052_ keymem.key_mem\[14\]\[56\]
+ _07963_ _08276_ sky130_fd_sc_hd__a221o_2
XFILLER_0_44_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16497_ VPWR VGND VGND VPWR _02657_ _02658_ _02656_ sky130_fd_sc_hd__nor2_2
XFILLER_0_31_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18236_ VPWR VGND VGND VPWR _04143_ _04140_ _04142_ sky130_fd_sc_hd__nand2_2
X_15448_ VPWR VGND _10909_ keymem.prev_key1_reg\[43\] keymem.prev_key1_reg\[11\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_217_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_127_387 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18167_ VGND VPWR _04080_ _03983_ _04079_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15379_ VGND VPWR VGND VPWR _10629_ _10608_ _10535_ _10515_ _10490_ _10840_ sky130_fd_sc_hd__o32a_2
XFILLER_0_142_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17118_ VGND VPWR VGND VPWR _03233_ _03231_ _03229_ _09534_ _03232_ _09514_ sky130_fd_sc_hd__a32o_2
XFILLER_0_40_333 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_111_86 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_223_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18098_ VPWR VGND VPWR VGND _04016_ block[99] _03980_ enc_block.block_w3_reg\[3\]
+ _04007_ _04017_ sky130_fd_sc_hd__a221o_2
XFILLER_0_1_920 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17049_ VPWR VGND VPWR VGND _03171_ _10086_ _03168_ _03169_ _03170_ _10096_ sky130_fd_sc_hd__o311a_2
XFILLER_0_187_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_141_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_964 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_110_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20060_ VGND VPWR VPWR VGND _05446_ _03075_ keymem.key_mem\[10\]\[52\] _05448_ sky130_fd_sc_hd__mux2_2
XFILLER_0_141_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Left_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_221_1270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_252_1208 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1339 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23750_ keymem.prev_key0_reg\[106\] clk _00247_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20962_ VPWR VGND keymem.key_mem\[7\]\[90\] _05928_ _05823_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_205_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22701_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[42\] _06790_ _06789_ _04939_ _02078_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_221_862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_152_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23681_ keymem.prev_key0_reg\[37\] clk _00178_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20893_ VGND VPWR VGND VPWR _05891_ keymem.key_mem_we _03119_ _05864_ _01197_ sky130_fd_sc_hd__a31o_2
XFILLER_0_221_873 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25420_ VGND VPWR VPWR VGND clk _01913_ reset_n keymem.key_mem\[1\]\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_152_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22632_ VGND VPWR VPWR VGND _06785_ keymem.key_mem\[0\]\[5\] _10194_ _06787_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_46_Left_314 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_113_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25351_ VGND VPWR VPWR VGND clk _01844_ reset_n keymem.key_mem\[2\]\[64\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_937 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22563_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[85\] _06754_ _06753_ _05008_ _01993_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_192_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24302_ VGND VPWR VPWR VGND clk _00795_ reset_n keymem.key_mem\[10\]\[39\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_1134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_118_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21514_ VGND VPWR _06220_ _06115_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25282_ VGND VPWR VPWR VGND clk _01775_ reset_n keymem.key_mem\[3\]\[123\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_17_Right_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22494_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[44\] _06737_ _06736_ _04943_ _01952_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_16_341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24233_ VGND VPWR VPWR VGND clk _00726_ reset_n keymem.key_mem\[11\]\[98\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21445_ VGND VPWR _06184_ _06115_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_9_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21376_ VGND VPWR VPWR VGND _06140_ _02786_ keymem.key_mem\[5\]\[28\] _06148_ sky130_fd_sc_hd__mux2_2
X_24164_ VGND VPWR VPWR VGND clk _00657_ reset_n keymem.key_mem\[11\]\[29\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_31_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1170 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_163_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23115_ VGND VPWR _02274_ _07036_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20327_ VGND VPWR _00933_ _05589_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24095_ VGND VPWR VPWR VGND clk _00588_ reset_n keymem.key_mem\[12\]\[88\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_222_1045 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_55_Left_323 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_60_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23046_ VGND VPWR VGND VPWR _02247_ _06994_ _06954_ keymem.prev_key1_reg\[70\] sky130_fd_sc_hd__o21a_2
XFILLER_0_120_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20258_ VGND VPWR _00900_ _05553_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_124_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_472 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_21_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20189_ VGND VPWR _05515_ _05387_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_26_Right_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_243_442 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24997_ VGND VPWR VPWR VGND clk _01490_ reset_n keymem.key_mem\[5\]\[94\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_263_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14750_ VGND VPWR VGND VPWR _09141_ _09136_ _09196_ _10216_ sky130_fd_sc_hd__a21o_2
X_23948_ VGND VPWR VPWR VGND clk _00441_ reset_n keymem.key_mem\[13\]\[69\] sky130_fd_sc_hd__dfrtp_2
X_11962_ VGND VPWR _07565_ _07564_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_192_1166 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_19_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13701_ VGND VPWR _09173_ _09172_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_170_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14681_ VPWR VGND VPWR VGND _09653_ _09970_ _09823_ _09225_ _10148_ sky130_fd_sc_hd__or4_2
XFILLER_0_54_1247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11893_ VGND VPWR result[113] _07510_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_64_Left_332 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23879_ VGND VPWR VPWR VGND clk _00372_ reset_n keymem.key_mem\[13\]\[0\] sky130_fd_sc_hd__dfrtp_2
X_16420_ VGND VPWR VGND VPWR _11345_ _11325_ _11306_ _11372_ _02582_ sky130_fd_sc_hd__a31o_2
XFILLER_0_131_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13632_ VGND VPWR VGND VPWR _09103_ _09095_ _09097_ _09100_ _09104_ sky130_fd_sc_hd__a31o_2
X_25618_ VGND VPWR VPWR VGND clk _02111_ reset_n keymem.key_mem\[0\]\[75\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_170_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_71_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_131_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16351_ VGND VPWR VGND VPWR _02514_ _02513_ _02512_ _02511_ _02510_ sky130_fd_sc_hd__and4_2
XFILLER_0_41_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13563_ VPWR VGND VPWR VGND _09014_ _09005_ _09034_ _09001_ _09035_ sky130_fd_sc_hd__or4_2
X_25549_ VGND VPWR VPWR VGND clk _02042_ reset_n keymem.key_mem\[0\]\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_55_948 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15302_ VPWR VGND VGND VPWR _10764_ _10472_ _10500_ sky130_fd_sc_hd__nand2_2
XFILLER_0_66_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12514_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[36\] _07588_ keymem.key_mem\[7\]\[36\]
+ _07610_ _08081_ sky130_fd_sc_hd__a22o_2
X_19070_ VPWR VGND keymem.key_mem\[13\]\[6\] _04888_ _04887_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16282_ VGND VPWR VGND VPWR _11239_ _11296_ _11253_ _11497_ _02446_ sky130_fd_sc_hd__o22a_2
X_13494_ enc_block.sword_ctr_reg\[1\] _08966_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[1\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_129_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18021_ VPWR VGND VGND VPWR _00000_ _03944_ _03945_ _00271_ sky130_fd_sc_hd__nor3_2
X_15233_ VPWR VGND VPWR VGND _10687_ _10695_ _10692_ _10681_ _10696_ sky130_fd_sc_hd__or4_2
XFILLER_0_212_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_23_812 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_124_346 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12445_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[30\] _07812_ keymem.key_mem\[4\]\[30\]
+ _07913_ _08018_ sky130_fd_sc_hd__a22o_2
X_15164_ VGND VPWR _10628_ _10469_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12376_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[24\] _07788_ keymem.key_mem\[1\]\[24\]
+ _07715_ _07955_ sky130_fd_sc_hd__a22o_2
XFILLER_0_209_1390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_889 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14115_ VGND VPWR VGND VPWR _09480_ _09559_ _09586_ _09563_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_181_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15095_ VGND VPWR _10559_ _10558_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19972_ VGND VPWR _00766_ _05401_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_142_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_266_545 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18923_ VPWR VGND VPWR VGND _04761_ _04664_ _04760_ enc_block.block_w2_reg\[17\]
+ _04709_ _00357_ sky130_fd_sc_hd__a221o_2
X_14046_ VPWR VGND VPWR VGND _09518_ key[0] _08935_ sky130_fd_sc_hd__or2_2
XFILLER_0_240_1178 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18854_ VPWR VGND VGND VPWR _04654_ _04700_ _04095_ sky130_fd_sc_hd__nor2_2
XFILLER_0_235_943 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_207_667 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_187_1_Right_788 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17805_ VPWR VGND VPWR VGND _03147_ _03799_ keymem.prev_key0_reg\[60\] _03788_ _00201_
+ sky130_fd_sc_hd__a22o_2
X_18785_ VGND VPWR _04637_ enc_block.block_w2_reg\[27\] _04636_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15997_ VPWR VGND VPWR VGND _11452_ _11450_ _11451_ sky130_fd_sc_hd__or2_2
XFILLER_0_261_250 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_235_998 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_234_486 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_37_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14948_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[9\] _09003_ _10412_ _09002_ _10390_
+ _10391_ sky130_fd_sc_hd__a32oi_2
X_17736_ VGND VPWR VPWR VGND _03723_ _02896_ keymem.prev_key0_reg\[35\] _03756_ sky130_fd_sc_hd__mux2_2
XFILLER_0_167_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14879_ _10342_ _10344_ _10340_ _10343_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_17667_ VGND VPWR VPWR VGND _03703_ _03707_ keymem.prev_key0_reg\[14\] _03708_ sky130_fd_sc_hd__mux2_2
XFILLER_0_15_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_253_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_207_Left_474 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19406_ VPWR VGND keymem.key_mem\[12\]\[3\] _05099_ _05095_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16618_ VGND VPWR _02774_ _02771_ _02773_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_17598_ VPWR VGND VGND VPWR _03656_ _03240_ _02823_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_53_Right_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_159_298 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16549_ VGND VPWR _02708_ _10278_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19337_ VPWR VGND keymem.key_mem_we _05052_ _03550_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_17_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_72_244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19268_ VGND VPWR _00456_ _05007_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_2_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1088 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_313 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_249_1170 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_801 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18219_ VGND VPWR _04127_ enc_block.block_w1_reg\[22\] enc_block.block_w0_reg\[30\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_182_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_823 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19199_ VPWR VGND keymem.key_mem\[13\]\[57\] _04966_ _04961_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_48_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_368 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21230_ VGND VPWR VPWR VGND _06065_ _03401_ keymem.key_mem\[6\]\[88\] _06070_ sky130_fd_sc_hd__mux2_2
XFILLER_0_40_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_216_Left_483 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21161_ VGND VPWR VPWR VGND _06029_ _03099_ keymem.key_mem\[6\]\[55\] _06034_ sky130_fd_sc_hd__mux2_2
XFILLER_0_1_750 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_145_1190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_62_Right_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20112_ VGND VPWR VPWR VGND _05469_ _03306_ keymem.key_mem\[10\]\[77\] _05475_ sky130_fd_sc_hd__mux2_2
X_21092_ VGND VPWR VPWR VGND _05996_ _02607_ keymem.key_mem\[6\]\[22\] _05998_ sky130_fd_sc_hd__mux2_2
XFILLER_0_0_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20043_ VGND VPWR VPWR VGND _05435_ _02998_ keymem.key_mem\[10\]\[44\] _05439_ sky130_fd_sc_hd__mux2_2
X_24920_ VGND VPWR VPWR VGND clk _01413_ reset_n keymem.key_mem\[5\]\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_256_1141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24851_ VGND VPWR VPWR VGND clk _01344_ reset_n keymem.key_mem\[6\]\[76\] sky130_fd_sc_hd__dfrtp_2
X_23802_ VGND VPWR VPWR VGND clk _00295_ reset_n enc_block.block_w0_reg\[21\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_648 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24782_ VGND VPWR VPWR VGND clk _01275_ reset_n keymem.key_mem\[6\]\[7\] sky130_fd_sc_hd__dfrtp_2
X_21994_ VGND VPWR VGND VPWR _06477_ keymem.key_mem_we _03150_ _06475_ _01712_ sky130_fd_sc_hd__a31o_2
XFILLER_0_94_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_225_Left_492 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23733_ keymem.prev_key0_reg\[89\] clk _00230_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20945_ VGND VPWR _01221_ _05919_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_152_1161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23664_ keymem.prev_key0_reg\[20\] clk _00161_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_48_230 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_95_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20876_ VGND VPWR _01189_ _05882_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_152_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25403_ VGND VPWR VPWR VGND clk _01896_ reset_n keymem.key_mem\[2\]\[116\] sky130_fd_sc_hd__dfrtp_2
X_22615_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[125\] _06756_ _03793_ _05085_ _02033_
+ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_115_2_Left_586 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_149_1_Right_750 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_948 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23595_ VGND VPWR VPWR VGND clk _00096_ reset_n keymem.key_mem\[14\]\[84\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_48_285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_447 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25334_ VGND VPWR VPWR VGND clk _01827_ reset_n keymem.key_mem\[2\]\[47\] sky130_fd_sc_hd__dfrtp_2
X_22546_ VGND VPWR _01981_ _06760_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_148_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_609 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_84_1_Left_351 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_84_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_267_1292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25265_ VGND VPWR VPWR VGND clk _01758_ reset_n keymem.key_mem\[3\]\[106\] sky130_fd_sc_hd__dfrtp_2
X_22477_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[32\] _06707_ _06706_ _04920_ _01940_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_121_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24216_ VGND VPWR VPWR VGND clk _00709_ reset_n keymem.key_mem\[11\]\[81\] sky130_fd_sc_hd__dfrtp_2
X_12230_ VGND VPWR VGND VPWR _07821_ _07665_ keymem.key_mem\[4\]\[12\] _07817_ _07820_
+ sky130_fd_sc_hd__a211o_2
X_21428_ VGND VPWR _01448_ _06175_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_241_1410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25196_ VGND VPWR VPWR VGND clk _01689_ reset_n keymem.key_mem\[3\]\[37\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_267_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24147_ VGND VPWR VPWR VGND clk _00640_ reset_n keymem.key_mem\[11\]\[12\] sky130_fd_sc_hd__dfrtp_2
X_12161_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[8\] _07610_ keymem.key_mem\[9\]\[8\]
+ _07593_ _07756_ sky130_fd_sc_hd__a22o_2
XFILLER_0_31_174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21359_ VGND VPWR VPWR VGND _06128_ _02479_ keymem.key_mem\[5\]\[20\] _06139_ sky130_fd_sc_hd__mux2_2
XFILLER_0_124_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_229_Right_98 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24078_ VGND VPWR VPWR VGND clk _00571_ reset_n keymem.key_mem\[12\]\[71\] sky130_fd_sc_hd__dfrtp_2
X_12092_ VGND VPWR _07690_ _07651_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_248_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15920_ VPWR VGND VGND VPWR _11376_ _11167_ _11265_ sky130_fd_sc_hd__nand2_2
XFILLER_0_25_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23029_ VGND VPWR VPWR VGND _06960_ _03192_ keymem.prev_key1_reg\[64\] _06984_ sky130_fd_sc_hd__mux2_2
XFILLER_0_263_537 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_21_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15851_ VPWR VGND VPWR VGND _11272_ _11229_ _11228_ _11225_ _11307_ sky130_fd_sc_hd__or4_2
XFILLER_0_102_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_95_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14802_ VPWR VGND VPWR VGND _10268_ keymem.prev_key0_reg\[6\] sky130_fd_sc_hd__inv_2
XFILLER_0_207_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15782_ VGND VPWR _11238_ _11237_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18570_ VPWR VGND _04444_ enc_block.block_w0_reg\[5\] enc_block.block_w3_reg\[13\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_12994_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[83\] _08137_ keymem.key_mem\[11\]\[83\]
+ _07809_ _08514_ sky130_fd_sc_hd__a22o_2
XFILLER_0_98_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14733_ VGND VPWR VPWR VGND _10000_ _10198_ _09834_ _10199_ sky130_fd_sc_hd__or3_2
X_17521_ VPWR VGND VGND VPWR _03589_ _02470_ _02471_ sky130_fd_sc_hd__nand2_2
XFILLER_0_203_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11945_ VGND VPWR VGND VPWR _07528_ _07548_ _07529_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_200_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17452_ VPWR VGND key[234] _03530_ _09522_ VPWR VGND sky130_fd_sc_hd__and2_2
X_14664_ VPWR VGND VGND VPWR _09564_ _09456_ _09396_ _09312_ _10131_ _10130_ sky130_fd_sc_hd__o221a_2
X_11876_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[9\] dec_new_block\[105\]
+ _07502_ sky130_fd_sc_hd__mux2_2
XFILLER_0_131_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16403_ VPWR VGND VGND VPWR _11268_ _11368_ _02564_ _02565_ sky130_fd_sc_hd__nor3_2
XFILLER_0_200_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13615_ VPWR VGND VGND VPWR _09086_ _09087_ _09051_ sky130_fd_sc_hd__nor2_2
XFILLER_0_71_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17383_ VPWR VGND VPWR VGND _03470_ key[97] _11543_ sky130_fd_sc_hd__or2_2
X_14595_ VPWR VGND VGND VPWR _09388_ _09375_ _10063_ _09373_ _09401_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_131_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_948 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19122_ VPWR VGND keymem.key_mem\[13\]\[29\] _04917_ _04915_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16334_ VGND VPWR _02497_ _02496_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_156_279 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_43_907 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13546_ VGND VPWR VPWR VGND _08963_ _09017_ _08957_ _09018_ sky130_fd_sc_hd__or3_2
XFILLER_0_32_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_767 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_166_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_469 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_55_778 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_124_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19053_ VGND VPWR _04877_ _04876_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16265_ VPWR VGND VPWR VGND _02425_ _02428_ _02429_ _11468_ _02423_ sky130_fd_sc_hd__or4b_2
XFILLER_0_36_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13477_ enc_block.sword_ctr_reg\[1\] _08949_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[2\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_15216_ VGND VPWR VGND VPWR _10539_ _10540_ _10530_ _10604_ _10679_ sky130_fd_sc_hd__o22a_2
X_18004_ VPWR VGND VPWR VGND _03645_ _03934_ keymem.prev_key0_reg\[124\] _03731_ _00265_
+ sky130_fd_sc_hd__a22o_2
X_12428_ VGND VPWR enc_block.round_key\[28\] _08002_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_2_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16196_ VGND VPWR VGND VPWR _02361_ _11494_ _11228_ _02359_ _02360_ sky130_fd_sc_hd__a211o_2
XFILLER_0_22_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15147_ VGND VPWR _10611_ _10610_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_11_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_24 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12359_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[22\] _07608_ keymem.key_mem\[9\]\[22\]
+ _07591_ _07940_ sky130_fd_sc_hd__a22o_2
XFILLER_0_199_1117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_103_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_267_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_77_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15078_ VGND VPWR VGND VPWR _10539_ _10538_ _10542_ _10541_ sky130_fd_sc_hd__a21oi_2
X_19955_ VGND VPWR _00758_ _05392_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_103_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14029_ _09407_ _09501_ _09364_ _09500_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_18906_ VGND VPWR _04746_ enc_block.block_w2_reg\[24\] _04745_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_177_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19886_ VGND VPWR _00727_ _05354_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_177_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18837_ VPWR VGND _04684_ enc_block.block_w0_reg\[15\] enc_block.block_w0_reg\[8\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_188_1_Right_789 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18768_ VPWR VGND _04622_ _04621_ enc_block.round_key\[34\] VPWR VGND sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_267_Right_136 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_136_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17719_ VPWR VGND VGND VPWR _03745_ _03746_ _03731_ sky130_fd_sc_hd__nor2_2
X_18699_ VPWR VGND VPWR VGND _04559_ _04550_ _04558_ enc_block.block_w1_reg\[27\]
+ _04328_ _00335_ sky130_fd_sc_hd__a221o_2
XFILLER_0_89_196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1166 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_77_347 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20730_ VGND VPWR _01124_ _05801_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_114_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_915 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_46_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_133_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_110_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20661_ VGND VPWR _01091_ _05765_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_50_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22400_ VGND VPWR _01904_ _06691_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_162_216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_11_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23380_ VPWR VGND _07254_ _07253_ enc_block.round_key\[17\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_20592_ VGND VPWR _01058_ _05729_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_18_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22331_ VGND VPWR _01871_ _06655_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_45_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_620 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_264_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25050_ VGND VPWR VPWR VGND clk _01543_ reset_n keymem.key_mem\[4\]\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_258 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22262_ VGND VPWR _01838_ _06619_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_5_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24001_ VGND VPWR VPWR VGND clk _00494_ reset_n keymem.key_mem\[13\]\[122\] sky130_fd_sc_hd__dfrtp_2
X_21213_ VGND VPWR VPWR VGND _06052_ _03329_ keymem.key_mem\[6\]\[80\] _06061_ sky130_fd_sc_hd__mux2_2
XFILLER_0_14_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22193_ VGND VPWR _01805_ _06583_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_44_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21144_ VGND VPWR VPWR VGND _06018_ _03024_ keymem.key_mem\[6\]\[47\] _06025_ sky130_fd_sc_hd__mux2_2
XFILLER_0_160_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_121_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_22_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_257_397 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21075_ VGND VPWR VPWR VGND _05983_ _11098_ keymem.key_mem\[6\]\[14\] _05989_ sky130_fd_sc_hd__mux2_2
XFILLER_0_195_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_226_740 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_22_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20026_ VGND VPWR VPWR VGND _05424_ _02913_ keymem.key_mem\[10\]\[36\] _05430_ sky130_fd_sc_hd__mux2_2
X_24903_ VGND VPWR VPWR VGND clk _01396_ reset_n keymem.key_mem\[5\]\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_201_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_784 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_233_Left_500 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24834_ VGND VPWR VPWR VGND clk _01327_ reset_n keymem.key_mem\[6\]\[59\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_234_Right_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_232_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24765_ VGND VPWR VPWR VGND clk _01258_ reset_n keymem.key_mem\[7\]\[118\] sky130_fd_sc_hd__dfrtp_2
X_21977_ VPWR VGND keymem.key_mem\[3\]\[53\] _06468_ _06439_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_95_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11730_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[0\] dec_new_block\[32\]
+ _07429_ sky130_fd_sc_hd__mux2_2
X_23716_ keymem.prev_key0_reg\[72\] clk _00213_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20928_ VGND VPWR VPWR VGND _05880_ _04989_ keymem.key_mem\[7\]\[74\] _05910_ sky130_fd_sc_hd__mux2_2
X_24696_ VGND VPWR VPWR VGND clk _01189_ reset_n keymem.key_mem\[7\]\[49\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_132_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_138_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11661_ VGND VPWR VGND VPWR _07395_ _07375_ _07394_ _07376_ enc_block.sword_ctr_inc
+ sky130_fd_sc_hd__and4_2
X_23647_ keymem.prev_key0_reg\[3\] clk _00144_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20859_ VGND VPWR _01181_ _05873_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13400_ VPWR VGND VPWR VGND _08879_ keymem.key_mem\[4\]\[123\] _07551_ keymem.key_mem\[2\]\[123\]
+ _07732_ _08880_ sky130_fd_sc_hd__a221o_2
X_14380_ VGND VPWR VGND VPWR _09838_ _09849_ _09850_ _09831_ _09845_ sky130_fd_sc_hd__nor4_2
XFILLER_0_36_244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23578_ VGND VPWR VPWR VGND clk _00079_ reset_n keymem.key_mem\[14\]\[67\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_91_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25317_ VGND VPWR VPWR VGND clk _01810_ reset_n keymem.key_mem\[2\]\[30\] sky130_fd_sc_hd__dfrtp_2
X_13331_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[116\] _07632_ keymem.key_mem\[11\]\[116\]
+ _07631_ _08818_ sky130_fd_sc_hd__a22o_2
X_22529_ VGND VPWR _01972_ _06752_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_51_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16050_ VGND VPWR VGND VPWR _11505_ _11503_ _11432_ _11341_ _11504_ sky130_fd_sc_hd__a211o_2
XFILLER_0_51_258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25248_ VGND VPWR VPWR VGND clk _01741_ reset_n keymem.key_mem\[3\]\[89\] sky130_fd_sc_hd__dfrtp_2
X_13262_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[109\] _07588_ keymem.key_mem\[3\]\[109\]
+ _07619_ _08756_ sky130_fd_sc_hd__a22o_2
XFILLER_0_121_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_243_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15001_ VPWR VGND VGND VPWR _10465_ _10463_ _10464_ sky130_fd_sc_hd__nand2_2
X_12213_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[11\] _07535_ _07804_ _07798_ _07805_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_32_472 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13193_ VGND VPWR VGND VPWR _08694_ _08096_ keymem.key_mem\[5\]\[102\] _08693_ _07573_
+ sky130_fd_sc_hd__a211o_2
X_25179_ VGND VPWR VPWR VGND clk _01672_ reset_n keymem.key_mem\[3\]\[20\] sky130_fd_sc_hd__dfrtp_2
X_12144_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[7\] _07595_ keymem.key_mem\[8\]\[7\]
+ _07654_ _07740_ sky130_fd_sc_hd__a22o_2
XFILLER_0_241_1284 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_678 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_206 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19740_ VGND VPWR VPWR VGND _05270_ keymem.key_mem\[11\]\[30\] _02839_ _05278_ sky130_fd_sc_hd__mux2_2
XFILLER_0_21_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16952_ VGND VPWR _03083_ _03082_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12075_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[3\] _07674_ keymem.key_mem\[12\]\[3\]
+ _07673_ _07675_ sky130_fd_sc_hd__a22o_2
XFILLER_0_198_1161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_159_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15903_ VGND VPWR VGND VPWR _11320_ _11313_ _11359_ _11238_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_21_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19671_ VGND VPWR _00627_ _05239_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_99_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16883_ VPWR VGND VGND VPWR _03020_ _10366_ _11144_ sky130_fd_sc_hd__nand2_2
X_18622_ VGND VPWR _04491_ _04488_ _04490_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15834_ VGND VPWR VGND VPWR _11290_ _11229_ _11289_ _11227_ _11288_ sky130_fd_sc_hd__and4_2
XFILLER_0_63_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18553_ VGND VPWR _04429_ _04426_ _04428_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15765_ VGND VPWR _11221_ _11216_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_86_100 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12977_ VGND VPWR VGND VPWR _07808_ keymem.key_mem\[12\]\[81\] _08496_ _08498_ _08499_
+ _08480_ sky130_fd_sc_hd__a2111o_2
X_17504_ VGND VPWR _00125_ _03574_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14716_ VPWR VGND VPWR VGND _09831_ _09996_ _09953_ _09696_ _10183_ sky130_fd_sc_hd__or4_2
X_11928_ VPWR VGND VGND VPWR _07531_ _07528_ _07529_ sky130_fd_sc_hd__nand2_2
X_18484_ VPWR VGND VPWR VGND _04367_ _04363_ _04365_ sky130_fd_sc_hd__or2_2
X_15696_ VGND VPWR VGND VPWR _10652_ _10552_ _11152_ keymem.prev_key1_reg\[112\] sky130_fd_sc_hd__a21oi_2
XFILLER_0_28_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_169_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_129_235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14647_ VGND VPWR VGND VPWR _09582_ _09480_ _10114_ _09486_ sky130_fd_sc_hd__a21oi_2
X_17435_ VPWR VGND VGND VPWR _03515_ key[232] _10278_ sky130_fd_sc_hd__nand2_2
X_11859_ VGND VPWR result[96] _07493_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_170_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14578_ VGND VPWR VPWR VGND _10043_ _10045_ _10041_ _10046_ sky130_fd_sc_hd__or3_2
X_17366_ VGND VPWR _09988_ keymem.prev_key0_reg\[95\] _03455_ _02847_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19105_ VGND VPWR VGND VPWR _04907_ keymem.key_mem_we _02550_ _04896_ _00393_ sky130_fd_sc_hd__a31o_2
X_13529_ VGND VPWR VGND VPWR _09001_ _08976_ _08975_ keymem.prev_key1_reg\[7\] _08969_
+ _08964_ sky130_fd_sc_hd__a32o_2
X_16317_ VGND VPWR VPWR VGND _11041_ keymem.key_mem\[14\]\[20\] _02480_ _02481_ sky130_fd_sc_hd__mux2_2
X_17297_ VGND VPWR VPWR VGND _03384_ keymem.key_mem\[14\]\[87\] _03393_ _03394_ sky130_fd_sc_hd__mux2_2
XFILLER_0_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1140 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19036_ VGND VPWR _04862_ enc_block.block_w3_reg\[21\] _04861_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_16248_ VGND VPWR VGND VPWR _10960_ _10948_ keymem.round_ctr_reg\[0\] _02412_ sky130_fd_sc_hd__a21o_2
XFILLER_0_152_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_67_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_623 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16179_ VPWR VGND _10861_ _02344_ _10892_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_242_1059 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_255_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19938_ VGND VPWR _00752_ _05381_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_195_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_278 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_208_751 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_78_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_103_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19869_ VGND VPWR _00719_ _05345_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_177_1267 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21900_ VGND VPWR VGND VPWR _06426_ keymem.key_mem_we _11547_ _06420_ _01669_ sky130_fd_sc_hd__a31o_2
XFILLER_0_78_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22880_ VGND VPWR VGND VPWR _06894_ _10145_ _03795_ _06884_ _10192_ sky130_fd_sc_hd__a211o_2
XFILLER_0_179_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21831_ VGND VPWR _01639_ _06387_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_253_1177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_218_1297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24550_ VGND VPWR VPWR VGND clk _01043_ reset_n keymem.key_mem\[8\]\[31\] sky130_fd_sc_hd__dfrtp_2
X_21762_ VGND VPWR _01606_ _06351_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23501_ VPWR VGND VPWR VGND _07360_ block[31] _03957_ enc_block.block_w3_reg\[31\]
+ _03952_ _07361_ sky130_fd_sc_hd__a221o_2
XFILLER_0_114_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20713_ VGND VPWR _01116_ _05792_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24481_ VGND VPWR VPWR VGND clk _00974_ reset_n keymem.key_mem\[9\]\[90\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_92_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21693_ VGND VPWR _01573_ _06315_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_11_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23432_ _07298_ _07300_ _07297_ _07299_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_50_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_149_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20644_ VGND VPWR _01083_ _05756_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_11_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_149_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23363_ VPWR VGND VPWR VGND _07238_ _04874_ _07237_ enc_block.block_w3_reg\[15\]
+ _07115_ _02320_ sky130_fd_sc_hd__a221o_2
XFILLER_0_6_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20575_ VGND VPWR _01050_ _05720_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_85_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25102_ VGND VPWR VPWR VGND clk _01595_ reset_n keymem.key_mem\[4\]\[71\] sky130_fd_sc_hd__dfrtp_2
X_22314_ VGND VPWR _01863_ _06646_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23294_ VPWR VGND _07176_ enc_block.block_w1_reg\[15\] enc_block.block_w1_reg\[8\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_103_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_85_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25033_ VGND VPWR VPWR VGND clk _01526_ reset_n keymem.key_mem\[4\]\[2\] sky130_fd_sc_hd__dfrtp_2
X_22245_ VGND VPWR _01830_ _06610_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_239_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22176_ VGND VPWR _01797_ _06574_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_125_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21127_ VGND VPWR VPWR VGND _06007_ _02945_ keymem.key_mem\[6\]\[39\] _06016_ sky130_fd_sc_hd__mux2_2
XFILLER_0_121_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21058_ VGND VPWR _01274_ _05979_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_156_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1367 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12900_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[73\] _08259_ _08429_ _08423_ _08430_
+ sky130_fd_sc_hd__o22a_2
X_20009_ VGND VPWR VPWR VGND _05413_ _02787_ keymem.key_mem\[10\]\[28\] _05421_ sky130_fd_sc_hd__mux2_2
X_13880_ VGND VPWR _09352_ _09351_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_96_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12831_ VGND VPWR enc_block.round_key\[66\] _08367_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24817_ VGND VPWR VPWR VGND clk _01310_ reset_n keymem.key_mem\[6\]\[42\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25797_ keymem.prev_key1_reg\[113\] clk _02290_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_198_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15550_ VPWR VGND VGND VPWR _10629_ _10583_ _10644_ _10513_ _11009_ _11008_ sky130_fd_sc_hd__o221a_2
X_12762_ VGND VPWR enc_block.round_key\[59\] _08305_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24748_ VGND VPWR VPWR VGND clk _01241_ reset_n keymem.key_mem\[7\]\[101\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_55_1172 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_57_818 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14501_ _09185_ _09970_ _09059_ _09666_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_11713_ VGND VPWR result[23] _07420_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_83_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_132_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15481_ VGND VPWR VPWR VGND _10772_ _10941_ _10940_ sky130_fd_sc_hd__and2b_2
X_24679_ VGND VPWR VPWR VGND clk _01172_ reset_n keymem.key_mem\[7\]\[32\] sky130_fd_sc_hd__dfrtp_2
X_12693_ VGND VPWR _08243_ _07746_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14432_ VGND VPWR VGND VPWR _09327_ _09565_ _09397_ _09487_ _09901_ sky130_fd_sc_hd__o22a_2
XFILLER_0_132_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17220_ VPWR VGND VPWR VGND _11155_ _11154_ key[208] _09866_ _03324_ sky130_fd_sc_hd__a22o_2
XFILLER_0_33_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11644_ VGND VPWR VGND VPWR _00007_ _07372_ enc_block.enc_ctrl_reg\[0\] _07377_ _07382_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_167_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_385 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_83_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17151_ VGND VPWR VPWR VGND _09517_ _10731_ keymem.prev_key0_reg\[73\] _03262_ sky130_fd_sc_hd__or3_2
XFILLER_0_167_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14363_ VGND VPWR VGND VPWR _09132_ _09174_ _09108_ _09087_ _09090_ _09833_ sky130_fd_sc_hd__o32a_2
XFILLER_0_68_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16102_ VGND VPWR VGND VPWR _11554_ _11553_ _11556_ _11555_ sky130_fd_sc_hd__a21oi_2
X_13314_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[114\] _08714_ _08802_ _08798_ _08803_
+ sky130_fd_sc_hd__o22a_2
X_17082_ VGND VPWR VGND VPWR _03200_ _09635_ _03201_ keylen sky130_fd_sc_hd__a21oi_2
X_14294_ VPWR VGND VPWR VGND _09762_ _09763_ _09764_ _09760_ _09761_ sky130_fd_sc_hd__or4b_2
XFILLER_0_247_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16033_ _11340_ _11488_ _11287_ _11417_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_33_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_243_1357 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_208_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13245_ VGND VPWR VGND VPWR _08741_ _08150_ keymem.key_mem\[3\]\[107\] _08738_ _08740_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_58_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13176_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[101\] _07894_ keymem.key_mem\[8\]\[101\]
+ _08211_ _08678_ sky130_fd_sc_hd__a22o_2
XFILLER_0_104_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1032 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_143_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12127_ VGND VPWR _07724_ _07595_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17984_ VGND VPWR VPWR VGND _03281_ key[246] keymem.prev_key1_reg\[118\] _03921_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_104_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_178_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19723_ VGND VPWR VPWR VGND _05259_ keymem.key_mem\[11\]\[22\] _02608_ _05269_ sky130_fd_sc_hd__mux2_2
XFILLER_0_100_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16935_ VGND VPWR _03068_ _03067_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12058_ VGND VPWR _07658_ _07598_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_174_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_849 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_75_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19654_ VGND VPWR VPWR VGND _05227_ _05073_ keymem.key_mem\[12\]\[119\] _05231_ sky130_fd_sc_hd__mux2_2
XFILLER_0_74_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16866_ VGND VPWR VPWR VGND _11034_ _03002_ _03005_ _02496_ _03004_ sky130_fd_sc_hd__o211a_2
XFILLER_0_254_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18605_ VPWR VGND _04476_ _04475_ enc_block.round_key\[81\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_75_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15817_ VGND VPWR _11273_ _11208_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19585_ VGND VPWR VPWR VGND _05183_ _05010_ keymem.key_mem\[12\]\[86\] _05195_ sky130_fd_sc_hd__mux2_2
XFILLER_0_215_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16797_ VGND VPWR VGND VPWR _09866_ key[167] _02942_ _02941_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_172_1153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_254_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18536_ VPWR VGND _04414_ _04413_ enc_block.round_key\[74\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_247_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15748_ VGND VPWR _11204_ _11203_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_115_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18467_ VGND VPWR _04351_ _03958_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15679_ VGND VPWR VPWR VGND _10885_ _11136_ _10811_ sky130_fd_sc_hd__and2b_2
XFILLER_0_23_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_74_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_8_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1508 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_12_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17418_ VGND VPWR _00113_ _03500_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_185_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_51_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18398_ VPWR VGND _04290_ _04289_ enc_block.round_key\[126\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_62_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_185_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17349_ VGND VPWR VGND VPWR _02793_ keymem.prev_key0_reg\[93\] _09517_ _03440_ sky130_fd_sc_hd__a21o_2
XFILLER_0_15_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_320 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_172_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_556 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_70_331 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20360_ VGND VPWR VPWR VGND _05602_ _03202_ keymem.key_mem\[9\]\[65\] _05607_ sky130_fd_sc_hd__mux2_2
XFILLER_0_226_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_130_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19019_ VGND VPWR _04847_ _04780_ _04846_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_183_1282 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_261_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20291_ VGND VPWR VPWR VGND _05569_ _02873_ keymem.key_mem\[9\]\[32\] _05571_ sky130_fd_sc_hd__mux2_2
XFILLER_0_2_174 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22030_ VGND VPWR _01729_ _06496_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_122_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_124_2_Left_595 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23981_ VGND VPWR VPWR VGND clk _00474_ reset_n keymem.key_mem\[13\]\[102\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_192_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_208_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25720_ keymem.prev_key1_reg\[36\] clk _02213_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_254_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22932_ VGND VPWR _06926_ _06880_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_93_1_Left_360 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_78_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25651_ VGND VPWR VPWR VGND clk _02144_ reset_n keymem.key_mem\[0\]\[108\] sky130_fd_sc_hd__dfrtp_2
X_22863_ VGND VPWR _06881_ _06880_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_35_1009 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_233_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24602_ VGND VPWR VPWR VGND clk _01095_ reset_n keymem.key_mem\[8\]\[83\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_937 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_167_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21814_ VGND VPWR VPWR VGND _06377_ _03538_ keymem.key_mem\[4\]\[107\] _06379_ sky130_fd_sc_hd__mux2_2
X_25582_ VGND VPWR VPWR VGND clk _02075_ reset_n keymem.key_mem\[0\]\[39\] sky130_fd_sc_hd__dfrtp_2
X_22794_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[97\] _06850_ _06849_ _05027_ _02133_
+ sky130_fd_sc_hd__a22o_2
X_24533_ VGND VPWR VPWR VGND clk _01026_ reset_n keymem.key_mem\[8\]\[14\] sky130_fd_sc_hd__dfrtp_2
X_21745_ VGND VPWR VGND VPWR _06259_ _03279_ _01598_ _06342_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_148_341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24464_ VGND VPWR VPWR VGND clk _00957_ reset_n keymem.key_mem\[9\]\[73\] sky130_fd_sc_hd__dfrtp_2
X_21676_ VGND VPWR _01565_ _06306_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_188_1171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23415_ VPWR VGND VGND VPWR _07285_ _07211_ _07284_ sky130_fd_sc_hd__nand2_2
X_20627_ VGND VPWR VPWR VGND _05747_ _03183_ keymem.key_mem\[8\]\[63\] _05748_ sky130_fd_sc_hd__mux2_2
XFILLER_0_190_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24395_ VGND VPWR VPWR VGND clk _00888_ reset_n keymem.key_mem\[9\]\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_61_342 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23346_ VGND VPWR _07223_ enc_block.block_w2_reg\[6\] _07222_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20558_ VGND VPWR _01042_ _05711_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_149_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_225_1054 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23277_ VPWR VGND VPWR VGND _07161_ _07157_ _07159_ sky130_fd_sc_hd__or2_2
X_20489_ VGND VPWR VPWR VGND _05534_ _03668_ keymem.key_mem\[9\]\[127\] _05674_ sky130_fd_sc_hd__mux2_2
X_13030_ VPWR VGND VPWR VGND _08546_ keymem.key_mem\[3\]\[86\] _08009_ keymem.key_mem\[2\]\[86\]
+ _07733_ _08547_ sky130_fd_sc_hd__a221o_2
X_25016_ VGND VPWR VPWR VGND clk _01509_ reset_n keymem.key_mem\[5\]\[113\] sky130_fd_sc_hd__dfrtp_2
X_22228_ VGND VPWR VPWR VGND _06600_ _02972_ keymem.key_mem\[2\]\[42\] _06602_ sky130_fd_sc_hd__mux2_2
XFILLER_0_30_795 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_266_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22159_ VGND VPWR _06565_ _06553_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_28_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14981_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[15\] _08989_ _10445_ _08983_ _10433_
+ _10434_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_234_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16720_ key[160] _02872_ keylen _10086_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_13932_ VGND VPWR _09404_ _09403_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_96_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13863_ VGND VPWR _09335_ _09334_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16651_ VGND VPWR VGND VPWR _02804_ _02803_ _02806_ _02805_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_212 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15602_ VGND VPWR VGND VPWR _10495_ _10437_ _11060_ _10489_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_57_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12814_ VPWR VGND VPWR VGND _08351_ keymem.key_mem\[14\]\[65\] _08003_ keymem.key_mem\[6\]\[65\]
+ _07771_ _08352_ sky130_fd_sc_hd__a221o_2
X_19370_ VGND VPWR _00491_ _05074_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_9_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13794_ VGND VPWR VGND VPWR _09266_ _09265_ _09264_ keymem.prev_key1_reg\[25\] _08989_
+ _08983_ sky130_fd_sc_hd__a32o_2
X_16582_ VPWR VGND VPWR VGND _02740_ key[154] _10286_ sky130_fd_sc_hd__or2_2
X_18321_ VPWR VGND VPWR VGND _04220_ block[118] _04213_ enc_block.block_w1_reg\[22\]
+ _04171_ _04221_ sky130_fd_sc_hd__a221o_2
XFILLER_0_201_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15533_ VPWR VGND VPWR VGND _10992_ _10936_ _10991_ sky130_fd_sc_hd__or2_2
X_12745_ VPWR VGND VPWR VGND _08289_ keymem.key_mem\[13\]\[58\] _07834_ keymem.key_mem\[14\]\[58\]
+ _08032_ _08290_ sky130_fd_sc_hd__a221o_2
XFILLER_0_38_840 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15464_ VGND VPWR VPWR VGND _10922_ _10923_ _10920_ _10924_ sky130_fd_sc_hd__or3_2
X_18252_ VPWR VGND _04158_ _04157_ enc_block.round_key\[112\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_56_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12676_ VPWR VGND VPWR VGND _08227_ keymem.key_mem\[13\]\[51\] _07730_ keymem.key_mem\[11\]\[51\]
+ _07902_ _08228_ sky130_fd_sc_hd__a221o_2
XFILLER_0_154_333 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14415_ VPWR VGND VGND VPWR _09487_ _09884_ _09456_ sky130_fd_sc_hd__nor2_2
X_17203_ VGND VPWR VGND VPWR _03308_ _11050_ _03309_ _11051_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_231_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_154_344 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11627_ VPWR VGND aes_core_ctrl_reg\[1\] _07368_ _07367_ VPWR VGND sky130_fd_sc_hd__and2_2
X_15395_ VPWR VGND VPWR VGND _10856_ _10485_ _10646_ sky130_fd_sc_hd__or2_2
X_18183_ VGND VPWR VGND VPWR _10814_ _10775_ _04073_ _04095_ sky130_fd_sc_hd__a21o_2
XFILLER_0_25_534 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_167_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14346_ VPWR VGND VPWR VGND _09810_ _09815_ _09812_ _09170_ _09816_ sky130_fd_sc_hd__or4_2
XFILLER_0_68_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17134_ VPWR VGND _10287_ _03247_ _10318_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_128_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_375 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17065_ VGND VPWR VPWR VGND _03185_ keymem.key_mem\[14\]\[63\] _03184_ _03186_ sky130_fd_sc_hd__mux2_2
X_14277_ VGND VPWR VGND VPWR _09564_ _09404_ _09747_ _09392_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16016_ VGND VPWR VGND VPWR _11379_ _11372_ _11298_ _11345_ _11471_ sky130_fd_sc_hd__o22a_2
X_13228_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[106\] _07872_ keymem.key_mem\[12\]\[106\]
+ _07620_ _08725_ sky130_fd_sc_hd__a22o_2
XFILLER_0_0_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_470 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_180_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_272 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1452 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13159_ VGND VPWR VGND VPWR _07778_ keymem.key_mem\[3\]\[99\] _08660_ _08662_ _08663_
+ _08599_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_197_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_104_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_225_827 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17967_ VGND VPWR _00253_ _03909_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_236_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19706_ VGND VPWR _00641_ _05260_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_139_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16918_ VGND VPWR VPWR VGND _10278_ key[178] keymem.prev_key1_reg\[50\] _03052_ sky130_fd_sc_hd__mux2_2
XFILLER_0_178_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_197_Right_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17898_ VGND VPWR VPWR VGND _03728_ _03862_ _03412_ _03863_ sky130_fd_sc_hd__or3_2
XFILLER_0_139_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19637_ VGND VPWR VPWR VGND _05216_ _05056_ keymem.key_mem\[12\]\[111\] _05222_ sky130_fd_sc_hd__mux2_2
X_16849_ VPWR VGND VPWR VGND _02989_ key[44] _10732_ sky130_fd_sc_hd__or2_2
XFILLER_0_251_178 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_75_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19568_ VGND VPWR VPWR VGND _05183_ _04997_ keymem.key_mem\[12\]\[78\] _05186_ sky130_fd_sc_hd__mux2_2
X_18519_ VGND VPWR VPWR VGND _04316_ enc_block.block_w1_reg\[8\] _04074_ _04399_ sky130_fd_sc_hd__mux2_2
XFILLER_0_8_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19499_ VGND VPWR VPWR VGND _05138_ _04947_ keymem.key_mem\[12\]\[46\] _05149_ sky130_fd_sc_hd__mux2_2
X_21530_ VGND VPWR _01497_ _06228_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_629 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_189_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21461_ VGND VPWR _06192_ _03227_ _01464_ _06114_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_7_266 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_12_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_320 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23200_ VPWR VGND _07091_ _07090_ enc_block.round_key\[0\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_248_1076 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20412_ VGND VPWR VPWR VGND _05627_ _03418_ keymem.key_mem\[9\]\[90\] _05634_ sky130_fd_sc_hd__mux2_2
XFILLER_0_86_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24180_ VGND VPWR VPWR VGND clk _00673_ reset_n keymem.key_mem\[11\]\[45\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21392_ VGND VPWR _01431_ _06156_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_146_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_515 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_70_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23131_ VGND VPWR VGND VPWR _03513_ _06928_ _03517_ _07046_ sky130_fd_sc_hd__a21o_2
X_20343_ VGND VPWR VPWR VGND _05591_ _03119_ keymem.key_mem\[9\]\[57\] _05598_ sky130_fd_sc_hd__mux2_2
XFILLER_0_47_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23062_ VGND VPWR VGND VPWR _02253_ _07004_ _06954_ keymem.prev_key1_reg\[76\] sky130_fd_sc_hd__o21a_2
XFILLER_0_45_1160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20274_ VGND VPWR VPWR VGND _05558_ _02689_ keymem.key_mem\[9\]\[24\] _05562_ sky130_fd_sc_hd__mux2_2
X_22013_ VGND VPWR VGND VPWR _06487_ keymem.key_mem_we _03235_ _06475_ _01721_ sky130_fd_sc_hd__a31o_2
XFILLER_0_216_827 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_227_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_259_1172 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_236_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23964_ VGND VPWR VPWR VGND clk _00457_ reset_n keymem.key_mem\[13\]\[85\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22915_ VGND VPWR VPWR VGND _06914_ _06913_ keymem.prev_key1_reg\[19\] _06915_ sky130_fd_sc_hd__mux2_2
X_25703_ keymem.prev_key1_reg\[19\] clk _02196_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_157_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23895_ VGND VPWR VPWR VGND clk _00388_ reset_n keymem.key_mem\[13\]\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25634_ VGND VPWR VPWR VGND clk _02127_ reset_n keymem.key_mem\[0\]\[91\] sky130_fd_sc_hd__dfrtp_2
X_22846_ VGND VPWR VGND VPWR keymem.rcon_logic.tmp_rcon\[0\] _06862_ keymem.rcon_logic.tmp_rcon\[7\]
+ _06863_ _02171_ sky130_fd_sc_hd__o22a_2
XFILLER_0_155_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25565_ VGND VPWR VPWR VGND clk _02058_ reset_n keymem.key_mem\[0\]\[22\] sky130_fd_sc_hd__dfrtp_2
X_22777_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[86\] _06850_ _06849_ _05010_ _02122_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_195_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12530_ VGND VPWR enc_block.round_key\[37\] _08095_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24516_ VGND VPWR VPWR VGND clk _01009_ reset_n keymem.key_mem\[9\]\[125\] sky130_fd_sc_hd__dfrtp_2
X_21728_ VGND VPWR VPWR VGND _06330_ _03209_ keymem.key_mem\[4\]\[66\] _06334_ sky130_fd_sc_hd__mux2_2
X_25496_ VGND VPWR VPWR VGND clk _01989_ reset_n keymem.key_mem\[1\]\[81\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_136_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24447_ VGND VPWR VPWR VGND clk _00940_ reset_n keymem.key_mem\[9\]\[56\] sky130_fd_sc_hd__dfrtp_2
X_12461_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[31\] _08032_ keymem.key_mem\[8\]\[31\]
+ _07929_ _08033_ sky130_fd_sc_hd__a22o_2
X_21659_ VGND VPWR VPWR VGND _06297_ _02883_ keymem.key_mem\[4\]\[33\] _06298_ sky130_fd_sc_hd__mux2_2
XFILLER_0_129_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14200_ VPWR VGND VGND VPWR _09196_ _09671_ _09071_ sky130_fd_sc_hd__nor2_2
XFILLER_0_168_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15180_ VGND VPWR _10644_ _10602_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_65_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12392_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[25\] _07619_ keymem.key_mem\[1\]\[25\]
+ _07969_ _07970_ sky130_fd_sc_hd__a22o_2
X_24378_ VGND VPWR VPWR VGND clk _00871_ reset_n keymem.key_mem\[10\]\[115\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_129_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_375 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_244_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14131_ VPWR VGND VGND VPWR _09408_ _09602_ _09375_ sky130_fd_sc_hd__nor2_2
XFILLER_0_209_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_846 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23329_ VPWR VGND VPWR VGND _07207_ block[12] _04837_ enc_block.block_w1_reg\[12\]
+ _04504_ _07208_ sky130_fd_sc_hd__a221o_2
XFILLER_0_65_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_210_Right_79 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14062_ VGND VPWR _09534_ _09533_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_39_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13013_ VGND VPWR enc_block.round_key\[84\] _08531_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18870_ VPWR VGND VGND VPWR _04713_ _04714_ _04478_ sky130_fd_sc_hd__nor2_2
XFILLER_0_123_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17821_ VGND VPWR _00207_ _03809_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_146_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17752_ VGND VPWR _00182_ _03765_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14964_ VPWR VGND VPWR VGND _10428_ enc_block.block_w0_reg\[14\] _09273_ sky130_fd_sc_hd__or2_2
XFILLER_0_262_977 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_136_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16703_ VGND VPWR _02856_ keymem.prev_key1_reg\[31\] keymem.prev_key1_reg\[63\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
X_13915_ VGND VPWR VPWR VGND _09304_ _09300_ _09297_ _09387_ sky130_fd_sc_hd__or3_2
XFILLER_0_251_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17683_ VGND VPWR _00160_ _03718_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_199_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1053 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14895_ VGND VPWR _10360_ _07386_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_255_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19422_ VGND VPWR VGND VPWR _05107_ keymem.key_mem_we _10836_ _05093_ _00510_ sky130_fd_sc_hd__a31o_2
XFILLER_0_18_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16634_ VGND VPWR VGND VPWR _02536_ _11301_ keymem.rcon_logic.tmp_rcon\[6\] _02789_
+ sky130_fd_sc_hd__a21o_2
X_13846_ VPWR VGND VPWR VGND _09299_ _09317_ _09315_ _09254_ _09318_ sky130_fd_sc_hd__or4_2
XFILLER_0_71_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_212_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19353_ VGND VPWR VPWR VGND _05046_ _05062_ keymem.key_mem\[13\]\[114\] _05063_ sky130_fd_sc_hd__mux2_2
X_13777_ VGND VPWR VGND VPWR _09249_ enc_block.block_w2_reg\[27\] enc_block.sword_ctr_reg\[1\]
+ enc_block.sword_ctr_reg\[0\] sky130_fd_sc_hd__and3b_2
X_16565_ VGND VPWR _02723_ _09543_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_146_108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18304_ VPWR VGND VPWR VGND _04205_ enc_block.block_w2_reg\[12\] enc_block.block_w2_reg\[13\]
+ sky130_fd_sc_hd__or2_2
XFILLER_0_70_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_127_311 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15516_ VGND VPWR VGND VPWR _08930_ key[140] _10975_ _10976_ sky130_fd_sc_hd__a21o_2
XFILLER_0_29_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19284_ VGND VPWR VGND VPWR _05017_ keymem.key_mem_we _03418_ _04999_ _00462_ sky130_fd_sc_hd__a31o_2
X_12728_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[56\] _07674_ keymem.key_mem\[1\]\[56\]
+ _07855_ _08275_ sky130_fd_sc_hd__a22o_2
XFILLER_0_112_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16496_ VGND VPWR VPWR VGND _09730_ _02650_ key[151] _02657_ sky130_fd_sc_hd__mux2_2
XFILLER_0_249_1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18235_ VGND VPWR _04142_ enc_block.block_w3_reg\[6\] _04141_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15447_ VPWR VGND VGND VPWR _10907_ _10908_ _10906_ sky130_fd_sc_hd__nor2_2
X_12659_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[50\] _07894_ keymem.key_mem\[8\]\[50\]
+ _08211_ _08212_ sky130_fd_sc_hd__a22o_2
XFILLER_0_142_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_112_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18166_ VPWR VGND _04079_ enc_block.block_w2_reg\[15\] enc_block.block_w2_reg\[8\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_15378_ _09941_ _10839_ _09240_ _09981_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_20_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17117_ VGND VPWR VPWR VGND _10322_ _10143_ key[197] _03232_ sky130_fd_sc_hd__mux2_2
X_14329_ VGND VPWR VGND VPWR _09799_ _09106_ _09798_ _09797_ sky130_fd_sc_hd__o21a_2
X_18097_ _04014_ _04016_ _04008_ _04015_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_20_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_223_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_932 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_208_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17048_ VPWR VGND VPWR VGND _03170_ key[190] _10322_ sky130_fd_sc_hd__or2_2
XFILLER_0_187_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_223_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_110_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18999_ VPWR VGND VPWR VGND _04829_ _04788_ _04828_ enc_block.block_w2_reg\[25\]
+ _04613_ _00365_ sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_150_2_Right_222 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_252_487 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20961_ VGND VPWR _01229_ _05927_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22700_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[41\] _06790_ _06789_ _04937_ _02077_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23680_ keymem.prev_key0_reg\[36\] clk _00177_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_7_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20892_ VPWR VGND keymem.key_mem\[7\]\[57\] _05891_ _05886_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_220_351 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22631_ VGND VPWR _02040_ _06786_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_467 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_75_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25350_ VGND VPWR VPWR VGND clk _01843_ reset_n keymem.key_mem\[2\]\[63\] sky130_fd_sc_hd__dfrtp_2
X_22562_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[84\] _06754_ _06753_ _05006_ _01992_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_118_322 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_267_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24301_ VGND VPWR VPWR VGND clk _00794_ reset_n keymem.key_mem\[10\]\[38\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_145_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21513_ VGND VPWR _01489_ _06219_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25281_ VGND VPWR VPWR VGND clk _01774_ reset_n keymem.key_mem\[3\]\[122\] sky130_fd_sc_hd__dfrtp_2
X_22493_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[43\] _06737_ _06736_ _04941_ _01951_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_118_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24232_ VGND VPWR VPWR VGND clk _00725_ reset_n keymem.key_mem\[11\]\[97\] sky130_fd_sc_hd__dfrtp_2
X_21444_ VGND VPWR _01456_ _06183_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_32_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_90_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_32_835 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24163_ VGND VPWR VPWR VGND clk _00656_ reset_n keymem.key_mem\[11\]\[28\] sky130_fd_sc_hd__dfrtp_2
X_21375_ VGND VPWR _01423_ _06147_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_31_356 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23114_ VGND VPWR VPWR VGND _07032_ _03473_ keymem.prev_key1_reg\[97\] _07036_ sky130_fd_sc_hd__mux2_2
XFILLER_0_82_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20326_ VGND VPWR VPWR VGND _05580_ _03046_ keymem.key_mem\[9\]\[49\] _05589_ sky130_fd_sc_hd__mux2_2
X_24094_ VGND VPWR VPWR VGND clk _00587_ reset_n keymem.key_mem\[12\]\[87\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_31_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23045_ VGND VPWR VGND VPWR _06994_ _03242_ _03241_ _03244_ _06951_ sky130_fd_sc_hd__a211o_2
X_20257_ VGND VPWR VPWR VGND _05546_ _11447_ keymem.key_mem\[9\]\[16\] _05553_ sky130_fd_sc_hd__mux2_2
XFILLER_0_228_440 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_200_1311 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_247_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20188_ VGND VPWR _00869_ _05514_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24996_ VGND VPWR VPWR VGND clk _01489_ reset_n keymem.key_mem\[5\]\[93\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_119_1_Left_386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_118_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11961_ VGND VPWR _07564_ _07563_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_19_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23947_ VGND VPWR VPWR VGND clk _00440_ reset_n keymem.key_mem\[13\]\[68\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13700_ VGND VPWR VPWR VGND _09031_ _08971_ _09008_ _09172_ sky130_fd_sc_hd__or3_2
X_14680_ VGND VPWR _10147_ keymem.prev_key0_reg\[5\] _10146_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_233_1131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_19_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11892_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[17\] dec_new_block\[113\]
+ _07510_ sky130_fd_sc_hd__mux2_2
X_23878_ VGND VPWR VPWR VGND clk _00371_ reset_n enc_block.block_w2_reg\[31\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13631_ VGND VPWR _09103_ _09102_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25617_ VGND VPWR VPWR VGND clk _02110_ reset_n keymem.key_mem\[0\]\[74\] sky130_fd_sc_hd__dfrtp_2
X_22829_ VPWR VGND VGND VPWR _06861_ _07387_ keylen sky130_fd_sc_hd__nand2_2
XFILLER_0_170_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16350_ VGND VPWR VGND VPWR _11319_ _11329_ _11245_ _11399_ _02513_ sky130_fd_sc_hd__o22a_2
X_13562_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[5\] _08956_ _09034_ _08943_ _08987_
+ _08988_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_66_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25548_ VGND VPWR VPWR VGND clk _02041_ reset_n keymem.key_mem\[0\]\[5\] sky130_fd_sc_hd__dfrtp_2
X_15301_ VPWR VGND VGND VPWR _10455_ _10763_ _10627_ sky130_fd_sc_hd__nor2_2
XFILLER_0_48_990 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12513_ VGND VPWR VGND VPWR _07580_ keymem.key_mem\[12\]\[36\] _08076_ _08079_ _08080_
+ _07574_ sky130_fd_sc_hd__a2111o_2
X_16281_ VGND VPWR VGND VPWR _11332_ _11375_ _11296_ _11469_ _02445_ sky130_fd_sc_hd__o22a_2
XFILLER_0_136_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13493_ VPWR VGND VGND VPWR enc_block.block_w1_reg\[1\] enc_block.sword_ctr_reg\[0\]
+ _08965_ sky130_fd_sc_hd__or2b_2
X_25479_ VGND VPWR VPWR VGND clk _01972_ reset_n keymem.key_mem\[1\]\[64\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_81_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_149_2_Left_620 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18020_ enc_block.round\[1\] _03945_ enc_block.round\[2\] _03941_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__and3_2
X_15232_ VPWR VGND VPWR VGND _10693_ _10694_ _10598_ _10505_ _10695_ sky130_fd_sc_hd__or4_2
XFILLER_0_129_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12444_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[30\] _07845_ keymem.key_mem\[6\]\[30\]
+ _07657_ _08017_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15163_ VGND VPWR _10627_ _10485_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12375_ VPWR VGND VPWR VGND _07953_ keymem.key_mem\[10\]\[24\] _07786_ keymem.key_mem\[4\]\[24\]
+ _07552_ _07954_ sky130_fd_sc_hd__a221o_2
XFILLER_0_1_228 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14114_ VGND VPWR VGND VPWR _09563_ _09450_ _09585_ _09582_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_26_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1282 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15094_ VPWR VGND VPWR VGND _10457_ _10445_ _10430_ _10443_ _10558_ sky130_fd_sc_hd__or4_2
X_19971_ VGND VPWR VPWR VGND _05400_ _10836_ keymem.key_mem\[10\]\[10\] _05401_ sky130_fd_sc_hd__mux2_2
XFILLER_0_181_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18922_ VPWR VGND VGND VPWR _04654_ _04761_ _04169_ sky130_fd_sc_hd__nor2_2
X_14045_ VGND VPWR _09517_ _09516_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_66_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_248_Right_117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_1063 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18853_ VPWR VGND _04699_ _04698_ enc_block.round_key\[42\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_234_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17804_ VPWR VGND VGND VPWR _03798_ _03799_ _03731_ sky130_fd_sc_hd__nor2_2
XFILLER_0_206_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18784_ VGND VPWR _04636_ enc_block.block_w2_reg\[31\] enc_block.block_w0_reg\[12\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15996_ _10677_ _11451_ keymem.prev_key1_reg\[113\] _10728_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_206_167 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17735_ VGND VPWR _00175_ _03755_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_222_627 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_221_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14947_ VGND VPWR _10411_ _10410_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_76_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_47 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17666_ VGND VPWR VPWR VGND _03691_ key[142] keymem.prev_key1_reg\[14\] _03707_ sky130_fd_sc_hd__mux2_2
XFILLER_0_37_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14878_ VGND VPWR VGND VPWR _09684_ _09167_ _09156_ _09029_ _10343_ sky130_fd_sc_hd__o22a_2
XFILLER_0_159_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19405_ VGND VPWR VGND VPWR _05098_ keymem.key_mem_we _09862_ _05093_ _00502_ sky130_fd_sc_hd__a31o_2
X_16617_ VGND VPWR _02773_ keymem.prev_key0_reg\[28\] _02772_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_13829_ VPWR VGND VPWR VGND _09299_ _09246_ _09300_ _09297_ _09301_ sky130_fd_sc_hd__or4_2
XFILLER_0_57_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_253_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17597_ VGND VPWR _00137_ _03655_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_9_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19336_ VGND VPWR _00480_ _05051_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_31_1023 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16548_ VGND VPWR VPWR VGND _02705_ _02691_ _02707_ _09514_ _02706_ sky130_fd_sc_hd__o211a_2
XFILLER_0_18_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_122_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19267_ VGND VPWR VPWR VGND _04993_ _05006_ keymem.key_mem\[13\]\[84\] _05007_ sky130_fd_sc_hd__mux2_2
X_16479_ VGND VPWR _02639_ _02610_ _02640_ _02638_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_31_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_45_459 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18218_ VGND VPWR VGND VPWR _04124_ _03951_ _04126_ _00287_ sky130_fd_sc_hd__a21o_2
XFILLER_0_147_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19198_ VGND VPWR VGND VPWR _04965_ keymem.key_mem_we _03109_ _04924_ _00428_ sky130_fd_sc_hd__a31o_2
XFILLER_0_108_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18149_ VPWR VGND VPWR VGND _04063_ _04040_ _04061_ enc_block.block_w0_reg\[7\] _03976_
+ _00281_ sky130_fd_sc_hd__a221o_2
XFILLER_0_40_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_643 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_2_Left_541 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21160_ VGND VPWR _01322_ _06033_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20111_ VGND VPWR _00832_ _05474_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21091_ VGND VPWR _01289_ _05997_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20042_ VGND VPWR _00799_ _05438_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_258_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24850_ VGND VPWR VPWR VGND clk _01343_ reset_n keymem.key_mem\[6\]\[75\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_2_Right_223 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23801_ VGND VPWR VPWR VGND clk _00294_ reset_n enc_block.block_w0_reg\[20\] sky130_fd_sc_hd__dfrtp_2
X_24781_ VGND VPWR VPWR VGND clk _01274_ reset_n keymem.key_mem\[6\]\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21993_ VPWR VGND keymem.key_mem\[3\]\[60\] _06477_ _06469_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_55_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23732_ keymem.prev_key0_reg\[88\] clk _00229_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20944_ VGND VPWR VPWR VGND _05912_ _05002_ keymem.key_mem\[7\]\[81\] _05919_ sky130_fd_sc_hd__mux2_2
XFILLER_0_95_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23663_ keymem.prev_key0_reg\[19\] clk _00160_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20875_ VGND VPWR VPWR VGND _05880_ _04953_ keymem.key_mem\[7\]\[49\] _05882_ sky130_fd_sc_hd__mux2_2
XFILLER_0_220_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_776 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22614_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[124\] _06756_ _03793_ _05083_ _02032_
+ sky130_fd_sc_hd__a22o_2
X_25402_ VGND VPWR VPWR VGND clk _01895_ reset_n keymem.key_mem\[2\]\[115\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_152_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_927 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_53_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23594_ VGND VPWR VPWR VGND clk _00095_ reset_n keymem.key_mem\[14\]\[83\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_118_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25333_ VGND VPWR VPWR VGND clk _01826_ reset_n keymem.key_mem\[2\]\[46\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_48_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22545_ VGND VPWR VPWR VGND _06750_ keymem.key_mem\[1\]\[73\] _03268_ _06760_ sky130_fd_sc_hd__mux2_2
XFILLER_0_64_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_118_163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25264_ VGND VPWR VPWR VGND clk _01757_ reset_n keymem.key_mem\[3\]\[105\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_133_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22476_ VGND VPWR _01939_ _06732_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_126_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24215_ VGND VPWR VPWR VGND clk _00708_ reset_n keymem.key_mem\[11\]\[80\] sky130_fd_sc_hd__dfrtp_2
X_21427_ VGND VPWR VPWR VGND _06173_ _03075_ keymem.key_mem\[5\]\[52\] _06175_ sky130_fd_sc_hd__mux2_2
XFILLER_0_224_1108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25195_ VGND VPWR VPWR VGND clk _01688_ reset_n keymem.key_mem\[3\]\[36\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_121_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12160_ VGND VPWR VGND VPWR _07755_ _07721_ keymem.key_mem\[14\]\[8\] _07754_ _07574_
+ sky130_fd_sc_hd__a211o_2
X_24146_ VGND VPWR VPWR VGND clk _00639_ reset_n keymem.key_mem\[11\]\[11\] sky130_fd_sc_hd__dfrtp_2
X_21358_ VGND VPWR _01415_ _06138_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_206_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_838 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_163_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20309_ VGND VPWR _05580_ _05534_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24077_ VGND VPWR VPWR VGND clk _00570_ reset_n keymem.key_mem\[12\]\[70\] sky130_fd_sc_hd__dfrtp_2
X_12091_ VGND VPWR enc_block.round_key\[4\] _07689_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_124_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21289_ VGND VPWR VPWR VGND _06098_ _03592_ keymem.key_mem\[6\]\[116\] _06101_ sky130_fd_sc_hd__mux2_2
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23028_ VGND VPWR VPWR VGND _02240_ _03177_ _03182_ _06925_ _06983_ sky130_fd_sc_hd__o31a_2
XFILLER_0_21_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_198_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15850_ VGND VPWR _11306_ _11305_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_774 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1362 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_95_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14801_ VGND VPWR VGND VPWR _10264_ _10263_ _10265_ _10267_ sky130_fd_sc_hd__a21o_2
X_15781_ VPWR VGND VPWR VGND _11206_ _11208_ _11197_ _11225_ _11237_ sky130_fd_sc_hd__or4_2
XFILLER_0_98_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_207_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24979_ VGND VPWR VPWR VGND clk _01472_ reset_n keymem.key_mem\[5\]\[76\] sky130_fd_sc_hd__dfrtp_2
X_12993_ VGND VPWR enc_block.round_key\[82\] _08513_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_203_126 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_19_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17520_ VGND VPWR VPWR VGND _10366_ _03587_ key[116] _03588_ sky130_fd_sc_hd__mux2_2
X_14732_ VPWR VGND VPWR VGND _10197_ _10198_ _09073_ _10196_ sky130_fd_sc_hd__or3b_2
X_11944_ VGND VPWR _07547_ _07546_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_213_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17451_ VGND VPWR VPWR VGND _03029_ _03528_ key[106] _03529_ sky130_fd_sc_hd__mux2_2
X_11875_ VGND VPWR result[104] _07501_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14663_ VGND VPWR VGND VPWR _09415_ _09479_ _09576_ _09408_ _10130_ sky130_fd_sc_hd__o22a_2
XFILLER_0_200_833 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_905 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_156_214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16402_ VGND VPWR VGND VPWR _11270_ _11246_ _02564_ _11527_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_131_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13614_ VGND VPWR _09086_ _09065_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17382_ VGND VPWR VPWR VGND _09710_ _09711_ _09932_ _03469_ sky130_fd_sc_hd__or3_2
X_14594_ VGND VPWR VGND VPWR _10061_ _10062_ _09756_ _09466_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_131_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19121_ VGND VPWR VGND VPWR _04916_ keymem.key_mem_we _02787_ _04908_ _00400_ sky130_fd_sc_hd__a31o_2
XFILLER_0_27_437 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_746 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16333_ VGND VPWR _02496_ _07378_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13545_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[1\] _08956_ _09017_ _08943_ _08967_
+ _08968_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_109_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19052_ VPWR VGND VGND VPWR _07387_ keymem.round_ctr_reg\[1\] _09538_ _04876_ sky130_fd_sc_hd__nor3_2
XFILLER_0_14_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16264_ VGND VPWR VPWR VGND _11372_ _11253_ _02428_ _02427_ _02426_ sky130_fd_sc_hd__o211a_2
X_13476_ VGND VPWR _08948_ _08947_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_54_278 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18003_ VPWR VGND VGND VPWR _03933_ _03934_ _03729_ sky130_fd_sc_hd__nor2_2
X_15215_ VPWR VGND VGND VPWR _10504_ _10527_ _10678_ _10563_ _10612_ sky130_fd_sc_hd__o22ai_2
X_12427_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[28\] _07644_ _08001_ _07997_ _08002_
+ sky130_fd_sc_hd__o22a_2
X_16195_ VGND VPWR VPWR VGND _11338_ _11395_ _02360_ _11417_ _11224_ sky130_fd_sc_hd__o211a_2
XFILLER_0_207_1339 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_267_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15146_ VPWR VGND VPWR VGND _10424_ _10435_ _10444_ _10443_ _10610_ sky130_fd_sc_hd__or4_2
XFILLER_0_267_822 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12358_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[22\] _07621_ keymem.key_mem\[1\]\[22\]
+ _07799_ _07939_ sky130_fd_sc_hd__a22o_2
XFILLER_0_142_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_77_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15077_ VGND VPWR _10541_ _10540_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19954_ VGND VPWR VPWR VGND _05389_ _09862_ keymem.key_mem\[10\]\[2\] _05392_ sky130_fd_sc_hd__mux2_2
X_12289_ VGND VPWR VGND VPWR _07737_ keymem.key_mem\[1\]\[17\] _07871_ _07874_ _07875_
+ _07663_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_142_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14028_ VGND VPWR VGND VPWR _09362_ _09319_ _09447_ _09500_ sky130_fd_sc_hd__a21o_2
X_18905_ VGND VPWR _04745_ enc_block.block_w3_reg\[23\] enc_block.block_w1_reg\[0\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19885_ VGND VPWR VPWR VGND _05350_ keymem.key_mem\[11\]\[99\] _03485_ _05354_ sky130_fd_sc_hd__mux2_2
XFILLER_0_219_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_207_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18836_ VPWR VGND _04683_ _04603_ enc_block.block_w1_reg\[1\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_184_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_235_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_306 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18767_ VPWR VGND VPWR VGND _04620_ block[34] _04576_ enc_block.block_w1_reg\[2\]
+ _04543_ _04621_ sky130_fd_sc_hd__a221o_2
X_15979_ VGND VPWR VGND VPWR _11349_ _11434_ _11327_ _11306_ _11435_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_89_142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_250_766 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17718_ VGND VPWR VGND VPWR _03732_ keymem.prev_key1_reg\[28\] _03745_ _03733_ sky130_fd_sc_hd__a21oi_2
X_18698_ VPWR VGND VGND VPWR _04512_ _04559_ _04258_ sky130_fd_sc_hd__nor2_2
XFILLER_0_72_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_194_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_212_1012 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_153_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17649_ VGND VPWR _00149_ _03695_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_147_214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_50_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20660_ VGND VPWR VPWR VGND _05761_ _03321_ keymem.key_mem\[8\]\[79\] _05765_ sky130_fd_sc_hd__mux2_2
XFILLER_0_147_247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_212_1089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19319_ VGND VPWR VPWR VGND _05025_ _05039_ keymem.key_mem\[13\]\[103\] _05040_ sky130_fd_sc_hd__mux2_2
X_20591_ VGND VPWR VPWR VGND _05725_ _03015_ keymem.key_mem\[8\]\[46\] _05729_ sky130_fd_sc_hd__mux2_2
XFILLER_0_2_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_821 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_11_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22330_ VGND VPWR VPWR VGND _06647_ _03426_ keymem.key_mem\[2\]\[91\] _06655_ sky130_fd_sc_hd__mux2_2
XFILLER_0_115_122 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_84_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22261_ VGND VPWR VPWR VGND _06611_ _03129_ keymem.key_mem\[2\]\[58\] _06619_ sky130_fd_sc_hd__mux2_2
XFILLER_0_264_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_665 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24000_ VGND VPWR VPWR VGND clk _00493_ reset_n keymem.key_mem\[13\]\[121\] sky130_fd_sc_hd__dfrtp_2
X_21212_ VGND VPWR _01347_ _06060_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_13_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_822 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22192_ VGND VPWR VPWR VGND _06578_ _02720_ keymem.key_mem\[2\]\[25\] _06583_ sky130_fd_sc_hd__mux2_2
XFILLER_0_160_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21143_ VGND VPWR _01314_ _06024_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_121_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_258_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_245_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_160_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_1_Left_535 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_121_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21074_ VGND VPWR _01281_ _05988_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_195_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20025_ VGND VPWR _00791_ _05429_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24902_ VGND VPWR VPWR VGND clk _01395_ reset_n keymem.key_mem\[6\]\[127\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24833_ VGND VPWR VPWR VGND clk _01326_ reset_n keymem.key_mem\[6\]\[58\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_225_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_244_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_152_2_Right_224 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21976_ VGND VPWR _01704_ _06467_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24764_ VGND VPWR VPWR VGND clk _01257_ reset_n keymem.key_mem\[7\]\[117\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_234_1270 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_197_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20927_ VGND VPWR VGND VPWR _05909_ keymem.key_mem_we _03268_ _05893_ _01213_ sky130_fd_sc_hd__a31o_2
X_23715_ keymem.prev_key0_reg\[71\] clk _00212_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_95_134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24695_ VGND VPWR VPWR VGND clk _01188_ reset_n keymem.key_mem\[7\]\[48\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_171_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_214 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_132_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11660_ VPWR VGND VGND VPWR enc_block.enc_ctrl_reg\[2\] _07394_ enc_block.enc_ctrl_reg\[3\]
+ sky130_fd_sc_hd__nor2_2
X_23646_ keymem.prev_key0_reg\[2\] clk _00143_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20858_ VGND VPWR VPWR VGND _05867_ _04937_ keymem.key_mem\[7\]\[41\] _05873_ sky130_fd_sc_hd__mux2_2
XFILLER_0_138_247 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23577_ VGND VPWR VPWR VGND clk _00078_ reset_n keymem.key_mem\[14\]\[66\] sky130_fd_sc_hd__dfrtp_2
X_20789_ VGND VPWR VGND VPWR _05835_ keymem.key_mem_we _10747_ _05821_ _01149_ sky130_fd_sc_hd__a31o_2
X_13330_ VPWR VGND VPWR VGND _08816_ keymem.key_mem\[6\]\[116\] _07657_ keymem.key_mem\[2\]\[116\]
+ _07698_ _08817_ sky130_fd_sc_hd__a221o_2
XFILLER_0_36_267 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22528_ VGND VPWR VPWR VGND _06750_ keymem.key_mem\[1\]\[64\] _03194_ _06752_ sky130_fd_sc_hd__mux2_2
X_25316_ VGND VPWR VPWR VGND clk _01809_ reset_n keymem.key_mem\[2\]\[29\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_91_373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_18_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_33_941 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13261_ VGND VPWR VGND VPWR _07737_ keymem.key_mem\[1\]\[109\] _08752_ _08754_ _08755_
+ _07896_ sky130_fd_sc_hd__a2111o_2
X_25247_ VGND VPWR VPWR VGND clk _01740_ reset_n keymem.key_mem\[3\]\[88\] sky130_fd_sc_hd__dfrtp_2
X_22459_ VGND VPWR _01931_ _06723_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_27_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_963 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15000_ VGND VPWR _10464_ _10409_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12212_ VGND VPWR VGND VPWR _07804_ _07800_ keymem.key_mem\[1\]\[11\] _07801_ _07803_
+ sky130_fd_sc_hd__a211o_2
X_13192_ VGND VPWR VGND VPWR _08693_ _07958_ keymem.key_mem\[8\]\[102\] _08690_ _08692_
+ sky130_fd_sc_hd__a211o_2
X_25178_ VGND VPWR VPWR VGND clk _01671_ reset_n keymem.key_mem\[3\]\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24129_ VGND VPWR VPWR VGND clk _00622_ reset_n keymem.key_mem\[12\]\[122\] sky130_fd_sc_hd__dfrtp_2
X_12143_ VGND VPWR _07739_ _07639_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_102_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_206_1394 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16951_ VGND VPWR VGND VPWR _08930_ key[181] _03081_ _03082_ sky130_fd_sc_hd__a21o_2
X_12074_ VGND VPWR _07674_ _07560_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_25_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15902_ VGND VPWR VGND VPWR _11358_ _11292_ _11287_ _11357_ _11349_ _11356_ sky130_fd_sc_hd__a32o_2
X_19670_ VGND VPWR VPWR VGND _05091_ _05089_ keymem.key_mem\[12\]\[127\] _05239_ sky130_fd_sc_hd__mux2_2
X_16882_ VGND VPWR VPWR VGND _11107_ _03018_ _03017_ _03019_ sky130_fd_sc_hd__mux2_2
XFILLER_0_159_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_379 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_21_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18621_ VGND VPWR _04490_ _04331_ _04489_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15833_ VGND VPWR _11289_ _11207_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_56_1107 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_154_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18552_ VPWR VGND _04428_ _04427_ _04355_ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_204_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15764_ VPWR VGND VGND VPWR _11182_ _11205_ _11220_ _11219_ _11211_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_38_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12976_ VPWR VGND VPWR VGND _08497_ keymem.key_mem\[7\]\[81\] _07650_ keymem.key_mem\[9\]\[81\]
+ _07738_ _08498_ sky130_fd_sc_hd__a221o_2
XFILLER_0_235_1078 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17503_ VGND VPWR VPWR VGND _03534_ keymem.key_mem\[14\]\[113\] _03573_ _03574_ sky130_fd_sc_hd__mux2_2
X_14715_ VPWR VGND VPWR VGND _10175_ _10181_ _10178_ _10172_ _10182_ sky130_fd_sc_hd__or4_2
XFILLER_0_59_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18483_ VPWR VGND VGND VPWR _04366_ _04363_ _04365_ sky130_fd_sc_hd__nand2_2
X_11927_ VPWR VGND VPWR VGND _07530_ _07528_ _07529_ sky130_fd_sc_hd__or2_2
XFILLER_0_169_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15695_ VGND VPWR _11151_ _09543_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17434_ VPWR VGND VGND VPWR _10374_ _03514_ _10373_ sky130_fd_sc_hd__nor2_2
X_14646_ _09478_ _10113_ _09360_ _09364_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_74_318 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_28_724 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11858_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[0\] dec_new_block\[96\]
+ _07493_ sky130_fd_sc_hd__mux2_2
XFILLER_0_86_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17365_ VPWR VGND keymem.prev_key0_reg\[95\] _03454_ _02847_ VPWR VGND sky130_fd_sc_hd__and2_2
X_14577_ VGND VPWR _10044_ _09333_ _10045_ _09341_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_11789_ VGND VPWR result[61] _07458_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_3_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19104_ VPWR VGND keymem.key_mem\[13\]\[21\] _04907_ _04903_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_12_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16316_ VGND VPWR _02480_ _02479_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_15_418 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13528_ VPWR VGND VGND VPWR _08999_ _09000_ _08972_ sky130_fd_sc_hd__nor2_2
X_17296_ VGND VPWR _03393_ _03392_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_12_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19035_ VGND VPWR _04861_ enc_block.block_w3_reg\[22\] enc_block.block_w1_reg\[6\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_952 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16247_ VGND VPWR _00031_ _02411_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_112_103 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13459_ VPWR VGND _08931_ keymem.prev_key0_reg\[64\] keymem.prev_key0_reg\[32\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_152_272 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_109_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16178_ VGND VPWR VGND VPWR _02343_ _09722_ _02342_ key[19] sky130_fd_sc_hd__o21a_2
XFILLER_0_11_635 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15129_ VGND VPWR _10593_ _10592_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_259_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19937_ VGND VPWR VPWR VGND _05372_ keymem.key_mem\[11\]\[124\] _03647_ _05381_ sky130_fd_sc_hd__mux2_2
XFILLER_0_220_1369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_79_1_Right_680 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_195_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_128_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_133_1_Left_400 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19868_ VGND VPWR VPWR VGND _05339_ keymem.key_mem\[11\]\[91\] _03427_ _05345_ sky130_fd_sc_hd__mux2_2
XFILLER_0_138_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18819_ VPWR VGND _04668_ enc_block.block_w2_reg\[31\] enc_block.block_w3_reg\[23\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_74_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19799_ VGND VPWR VPWR VGND _05303_ keymem.key_mem\[11\]\[58\] _03130_ _05309_ sky130_fd_sc_hd__mux2_2
XFILLER_0_78_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_179_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_253_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21830_ VGND VPWR VPWR VGND _06377_ _03585_ keymem.key_mem\[4\]\[115\] _06387_ sky130_fd_sc_hd__mux2_2
XFILLER_0_223_777 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_223_788 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21761_ VGND VPWR VPWR VGND _06344_ _03346_ keymem.key_mem\[4\]\[82\] _06351_ sky130_fd_sc_hd__mux2_2
XFILLER_0_19_702 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23500_ _07358_ _07360_ _03981_ _07359_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_20712_ VGND VPWR VPWR VGND _05783_ _03518_ keymem.key_mem\[8\]\[104\] _05792_ sky130_fd_sc_hd__mux2_2
XFILLER_0_53_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24480_ VGND VPWR VPWR VGND clk _00973_ reset_n keymem.key_mem\[9\]\[89\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_114_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21692_ VGND VPWR VPWR VGND _06308_ _03046_ keymem.key_mem\[4\]\[49\] _06315_ sky130_fd_sc_hd__mux2_2
XFILLER_0_46_510 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23431_ VPWR VGND VPWR VGND _07299_ enc_block.block_w3_reg\[31\] enc_block.block_w1_reg\[14\]
+ sky130_fd_sc_hd__or2_2
XFILLER_0_92_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20643_ VGND VPWR VPWR VGND _05747_ _03251_ keymem.key_mem\[8\]\[71\] _05756_ sky130_fd_sc_hd__mux2_2
XFILLER_0_11_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23362_ VPWR VGND VGND VPWR _07192_ _07238_ _04137_ sky130_fd_sc_hd__nor2_2
XFILLER_0_85_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20574_ VGND VPWR VPWR VGND _05714_ _02934_ keymem.key_mem\[8\]\[38\] _05720_ sky130_fd_sc_hd__mux2_2
XFILLER_0_149_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_662 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22313_ VGND VPWR VPWR VGND _06634_ _03355_ keymem.key_mem\[2\]\[83\] _06646_ sky130_fd_sc_hd__mux2_2
X_25101_ VGND VPWR VPWR VGND clk _01594_ reset_n keymem.key_mem\[4\]\[70\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_150_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23293_ VGND VPWR _07175_ enc_block.block_w2_reg\[1\] _07098_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_128_1_Left_395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25032_ VGND VPWR VPWR VGND clk _01525_ reset_n keymem.key_mem\[4\]\[1\] sky130_fd_sc_hd__dfrtp_2
X_22244_ VGND VPWR VPWR VGND _06600_ _03056_ keymem.key_mem\[2\]\[50\] _06610_ sky130_fd_sc_hd__mux2_2
XFILLER_0_41_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1033 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22175_ VGND VPWR VPWR VGND _06565_ _11546_ keymem.key_mem\[2\]\[17\] _06574_ sky130_fd_sc_hd__mux2_2
XFILLER_0_2_890 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21126_ VGND VPWR _01306_ _06015_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_160_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21057_ VGND VPWR VPWR VGND _05972_ _10283_ keymem.key_mem\[6\]\[6\] _05979_ sky130_fd_sc_hd__mux2_2
XFILLER_0_255_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_156_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20008_ VGND VPWR _00783_ _05420_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_92_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12830_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[66\] _08259_ _08366_ _08360_ _08367_
+ sky130_fd_sc_hd__o22a_2
X_24816_ VGND VPWR VPWR VGND clk _01309_ reset_n keymem.key_mem\[6\]\[41\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_214_777 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25796_ keymem.prev_key1_reg\[112\] clk _02289_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_153_2_Right_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_119_1174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12761_ VGND VPWR VGND VPWR _07793_ keymem.key_mem\[0\]\[59\] _08304_ _08300_ _08298_
+ _08305_ sky130_fd_sc_hd__o32a_2
X_24747_ VGND VPWR VPWR VGND clk _01240_ reset_n keymem.key_mem\[7\]\[100\] sky130_fd_sc_hd__dfrtp_2
X_21959_ VGND VPWR _01696_ _06458_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_201_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14500_ VPWR VGND VGND VPWR _09100_ _09969_ _09149_ sky130_fd_sc_hd__nor2_2
X_11712_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[23\] dec_new_block\[23\]
+ _07420_ sky130_fd_sc_hd__mux2_2
X_15480_ VGND VPWR VGND VPWR _10603_ _10568_ _10594_ _10478_ _10514_ _10940_ sky130_fd_sc_hd__o32a_2
X_12692_ VPWR VGND VPWR VGND _08241_ keymem.key_mem\[5\]\[53\] _07811_ keymem.key_mem\[9\]\[53\]
+ _07738_ _08242_ sky130_fd_sc_hd__a221o_2
XFILLER_0_132_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24678_ VGND VPWR VPWR VGND clk _01171_ reset_n keymem.key_mem\[7\]\[31\] sky130_fd_sc_hd__dfrtp_2
X_14431_ VGND VPWR VGND VPWR _09268_ _09330_ _09426_ _09582_ _09248_ _09900_ sky130_fd_sc_hd__o32a_2
X_11643_ VPWR VGND VPWR VGND _07382_ _07381_ sky130_fd_sc_hd__inv_2
X_23629_ VGND VPWR VPWR VGND clk _00130_ reset_n keymem.key_mem\[14\]\[118\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_167_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17150_ VPWR VGND VPWR VGND _10740_ _10739_ key[201] _09866_ _03261_ sky130_fd_sc_hd__a22o_2
XFILLER_0_37_587 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14362_ VGND VPWR VGND VPWR _09056_ _09687_ _09095_ _09100_ _09832_ sky130_fd_sc_hd__a31o_2
XFILLER_0_167_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16101_ VPWR VGND VPWR VGND _11555_ keymem.prev_key1_reg\[82\] sky130_fd_sc_hd__inv_2
X_13313_ VGND VPWR VGND VPWR _08802_ _07839_ keymem.key_mem\[11\]\[114\] _08799_ _08801_
+ sky130_fd_sc_hd__a211o_2
X_14293_ VGND VPWR VPWR VGND _09310_ _09407_ _09362_ _09763_ sky130_fd_sc_hd__or3_2
X_17081_ VPWR VGND VGND VPWR _03200_ key[193] _03077_ sky130_fd_sc_hd__nand2_2
XFILLER_0_40_719 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16032_ _11477_ _11487_ _11223_ _11426_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_13244_ VPWR VGND VPWR VGND _08739_ keymem.key_mem\[13\]\[107\] _08125_ keymem.key_mem\[2\]\[107\]
+ _07647_ _08740_ sky130_fd_sc_hd__a221o_2
XFILLER_0_126_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_630 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13175_ VGND VPWR enc_block.round_key\[100\] _08677_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_21_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12126_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[6\] _07668_ keymem.key_mem\[12\]\[6\]
+ _07722_ _07723_ sky130_fd_sc_hd__a22o_2
XFILLER_0_209_538 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17983_ VGND VPWR _00258_ _03920_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_100_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19722_ VGND VPWR _00649_ _05268_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_40_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16934_ VGND VPWR VGND VPWR _03066_ key[179] _03067_ _11151_ sky130_fd_sc_hd__a21bo_2
X_12057_ VGND VPWR _07657_ _07656_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_178_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_74_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19653_ VGND VPWR _00618_ _05230_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16865_ VGND VPWR VGND VPWR _11033_ _11032_ _03003_ _03004_ sky130_fd_sc_hd__a21o_2
XFILLER_0_217_593 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_204_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18604_ VPWR VGND VPWR VGND _04474_ block[81] _04330_ enc_block.block_w2_reg\[17\]
+ _04425_ _04475_ sky130_fd_sc_hd__a221o_2
X_15816_ VGND VPWR _11272_ _11206_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_254_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19584_ VGND VPWR _00585_ _05194_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16796_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[71\] keymem.prev_key1_reg\[39\]
+ _02941_ _02940_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_99_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_149_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18535_ VPWR VGND VPWR VGND _04412_ block[74] _04330_ enc_block.block_w3_reg\[10\]
+ _04276_ _04413_ sky130_fd_sc_hd__a221o_2
XFILLER_0_181_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15747_ VPWR VGND VPWR VGND _11192_ _11202_ _11197_ _11187_ _11203_ sky130_fd_sc_hd__or4_2
X_12959_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[79\] _07632_ keymem.key_mem\[9\]\[79\]
+ _07612_ _08483_ sky130_fd_sc_hd__a22o_2
XFILLER_0_59_156 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_142_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_252_Left_519 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18466_ VGND VPWR _04350_ _04019_ _00311_ _04317_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_15678_ VGND VPWR VGND VPWR _11135_ _11134_ _11129_ _11126_ _11125_ sky130_fd_sc_hd__and4_2
XFILLER_0_47_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_111_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_54 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_115_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_150_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17417_ VGND VPWR VPWR VGND _03467_ keymem.key_mem\[14\]\[101\] _03499_ _03500_ sky130_fd_sc_hd__mux2_2
X_14629_ VPWR VGND VPWR VGND _10097_ _10086_ _10089_ _10090_ _10095_ _10096_ sky130_fd_sc_hd__o311a_2
XFILLER_0_8_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18397_ VPWR VGND VPWR VGND _04288_ block[126] _04213_ enc_block.block_w0_reg\[30\]
+ _04276_ _04289_ sky130_fd_sc_hd__a221o_2
XFILLER_0_111_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_185_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17348_ VPWR VGND VGND VPWR _02793_ _03439_ keymem.prev_key0_reg\[93\] sky130_fd_sc_hd__nor2_2
XFILLER_0_12_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_209_1209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_172_356 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_185_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_265_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_248 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_70_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17279_ VGND VPWR keymem.prev_key0_reg\[86\] _02588_ _03377_ _02589_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_130_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19018_ VPWR VGND _04846_ enc_block.block_w1_reg\[4\] enc_block.block_w3_reg\[20\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_3_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20290_ VGND VPWR _00915_ _05570_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_11_410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_933 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_259_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_261_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_100_106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_261_Left_528 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_122_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1310 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_139_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_227_346 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_47_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23980_ VGND VPWR VPWR VGND clk _00473_ reset_n keymem.key_mem\[13\]\[101\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_192_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22931_ VGND VPWR _06925_ _06924_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_78_1162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_155_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_233_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_78_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25650_ VGND VPWR VPWR VGND clk _02143_ reset_n keymem.key_mem\[0\]\[107\] sky130_fd_sc_hd__dfrtp_2
X_22862_ VGND VPWR _06880_ _06877_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_64_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24601_ VGND VPWR VPWR VGND clk _01094_ reset_n keymem.key_mem\[8\]\[82\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_233_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21813_ VGND VPWR _01630_ _06378_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_196_949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22793_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[96\] _06850_ _06849_ _05024_ _02132_
+ sky130_fd_sc_hd__a22o_2
X_25581_ VGND VPWR VPWR VGND clk _02074_ reset_n keymem.key_mem\[0\]\[38\] sky130_fd_sc_hd__dfrtp_2
X_21744_ VPWR VGND VGND VPWR _06259_ _06342_ keymem.key_mem\[4\]\[74\] sky130_fd_sc_hd__nor2_2
X_24532_ VGND VPWR VPWR VGND clk _01025_ reset_n keymem.key_mem\[8\]\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_65_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21675_ VGND VPWR VPWR VGND _06297_ _02964_ keymem.key_mem\[4\]\[41\] _06306_ sky130_fd_sc_hd__mux2_2
X_24463_ VGND VPWR VPWR VGND clk _00956_ reset_n keymem.key_mem\[9\]\[72\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_148_386 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23414_ VGND VPWR _07284_ enc_block.block_w1_reg\[13\] _07283_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20626_ VGND VPWR _05747_ _05679_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_34_513 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24394_ VGND VPWR VPWR VGND clk _00887_ reset_n keymem.key_mem\[9\]\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_149_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23345_ VGND VPWR _07222_ enc_block.block_w2_reg\[5\] enc_block.block_w1_reg\[13\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20557_ VGND VPWR VPWR VGND _05703_ _02838_ keymem.key_mem\[8\]\[30\] _05711_ sky130_fd_sc_hd__mux2_2
XFILLER_0_61_354 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_62_899 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23276_ VPWR VGND VGND VPWR _07160_ _07157_ _07159_ sky130_fd_sc_hd__nand2_2
XFILLER_0_264_1093 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_85_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20488_ VGND VPWR _01010_ _05673_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22227_ VGND VPWR _01821_ _06601_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25015_ VGND VPWR VPWR VGND clk _01508_ reset_n keymem.key_mem\[5\]\[112\] sky130_fd_sc_hd__dfrtp_2
X_22158_ VGND VPWR _01789_ _06564_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21109_ VGND VPWR _01298_ _06006_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14980_ VGND VPWR VGND VPWR _10444_ _10428_ _10427_ keymem.prev_key1_reg\[14\] _09003_
+ _09002_ sky130_fd_sc_hd__a32o_2
X_22089_ VGND VPWR _06527_ _06402_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_22_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13931_ VGND VPWR _09403_ _09402_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_199_710 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_96_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16650_ VGND VPWR _02805_ keymem.prev_key1_reg\[29\] keymem.prev_key1_reg\[61\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
X_13862_ VPWR VGND VPWR VGND _09280_ _09291_ _09321_ _09275_ _09334_ sky130_fd_sc_hd__or4_2
XFILLER_0_44_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_168 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_57_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_138_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15601_ VGND VPWR VGND VPWR _10495_ _10476_ _11059_ _10602_ sky130_fd_sc_hd__a21oi_2
X_12813_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[65\] _07812_ keymem.key_mem\[4\]\[65\]
+ _07636_ _08351_ sky130_fd_sc_hd__a22o_2
XFILLER_0_241_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16581_ VGND VPWR VGND VPWR _02736_ _02735_ _02739_ _02737_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_158_117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13793_ VPWR VGND VPWR VGND _09265_ enc_block.block_w0_reg\[25\] _08952_ sky130_fd_sc_hd__or2_2
X_25779_ keymem.prev_key1_reg\[95\] clk _02272_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_154_2_Right_226 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_74_1582 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_198_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18320_ VGND VPWR VGND VPWR _04220_ _03982_ _04219_ _04218_ sky130_fd_sc_hd__o21a_2
X_15532_ VPWR VGND VPWR VGND _10989_ _10990_ _10991_ _10721_ _10988_ sky130_fd_sc_hd__or4b_2
X_12744_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[58\] _07659_ keymem.key_mem\[1\]\[58\]
+ _07714_ _08289_ sky130_fd_sc_hd__a22o_2
XFILLER_0_139_353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18251_ VPWR VGND VPWR VGND _04156_ block[112] _04076_ enc_block.block_w1_reg\[16\]
+ _04007_ _04157_ sky130_fd_sc_hd__a221o_2
XFILLER_0_132_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15463_ VGND VPWR VPWR VGND _10781_ _10782_ _10542_ _10923_ sky130_fd_sc_hd__or3_2
XFILLER_0_166_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12675_ VPWR VGND VPWR VGND keymem.key_mem\[8\]\[51\] _07752_ keymem.key_mem\[1\]\[51\]
+ _07855_ _08227_ sky130_fd_sc_hd__a22o_2
X_17202_ VPWR VGND VGND VPWR _03308_ key[206] _10278_ sky130_fd_sc_hd__nand2_2
X_14414_ VPWR VGND VGND VPWR _09875_ _09878_ _09882_ _09883_ sky130_fd_sc_hd__nor3_2
X_18182_ VPWR VGND _04094_ _04093_ enc_block.round_key\[106\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_11626_ VGND VPWR VPWR VGND encdec enc_block.ready dec_ready _07367_ sky130_fd_sc_hd__mux2_2
X_15394_ VPWR VGND VPWR VGND _10753_ _10854_ _10851_ _10640_ _10855_ sky130_fd_sc_hd__or4_2
XFILLER_0_68_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_167_1245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_114_209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_128_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17133_ VGND VPWR _00082_ _03246_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_167_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14345_ VGND VPWR VGND VPWR _09815_ _09672_ _09181_ _09813_ _09814_ sky130_fd_sc_hd__a211o_2
XFILLER_0_107_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17064_ VGND VPWR _03185_ _09863_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14276_ VPWR VGND VGND VPWR _09359_ _09427_ _09741_ _09745_ _09746_ sky130_fd_sc_hd__and4b_2
XFILLER_0_122_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_243_1166 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_204_1117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16015_ VGND VPWR VGND VPWR _11345_ _11466_ _11296_ _11469_ _11470_ sky130_fd_sc_hd__o22a_2
XFILLER_0_21_741 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13227_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[106\] _07919_ keymem.key_mem\[1\]\[106\]
+ _07715_ _08724_ sky130_fd_sc_hd__a22o_2
XFILLER_0_100_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13158_ VPWR VGND VPWR VGND _08661_ keymem.key_mem\[5\]\[99\] _07811_ keymem.key_mem\[7\]\[99\]
+ _07609_ _08662_ sky130_fd_sc_hd__a221o_2
XFILLER_0_20_284 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_430 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_209_346 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12109_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[5\] _07674_ keymem.key_mem\[1\]\[5\]
+ _07557_ _07707_ sky130_fd_sc_hd__a22o_2
X_17966_ VGND VPWR VPWR VGND _03896_ _03908_ keymem.prev_key0_reg\[112\] _03909_ sky130_fd_sc_hd__mux2_2
X_13089_ VGND VPWR VGND VPWR _07908_ keymem.key_mem\[6\]\[92\] _08596_ _08598_ _08600_
+ _08599_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_40_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_237_699 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16917_ VPWR VGND VGND VPWR _11557_ _03051_ _11556_ sky130_fd_sc_hd__nor2_2
X_19705_ VGND VPWR VPWR VGND _05259_ keymem.key_mem\[11\]\[13\] _11040_ _05260_ sky130_fd_sc_hd__mux2_2
XFILLER_0_79_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17897_ VGND VPWR VGND VPWR _03737_ keymem.prev_key1_reg\[90\] _03862_ _03738_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_139_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_850 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_189_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_75_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16848_ VPWR VGND VPWR VGND _02988_ _10915_ sky130_fd_sc_hd__inv_2
XFILLER_0_219_1371 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19636_ VGND VPWR _00610_ _05221_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_75_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19567_ VGND VPWR _00577_ _05185_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16779_ VGND VPWR _00049_ _02925_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18518_ VPWR VGND _04398_ _04397_ enc_block.round_key\[72\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_19498_ VGND VPWR _00545_ _05148_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_8_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18449_ VPWR VGND VGND VPWR _04335_ _04331_ _04333_ sky130_fd_sc_hd__nand2_2
XFILLER_0_115_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_735 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_111_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21460_ VPWR VGND VGND VPWR _06192_ keymem.key_mem\[5\]\[68\] _06114_ sky130_fd_sc_hd__nand2_2
XFILLER_0_86_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_546 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20411_ VGND VPWR _00973_ _05633_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_146_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21391_ VGND VPWR VPWR VGND _06151_ _02903_ keymem.key_mem\[5\]\[35\] _06156_ sky130_fd_sc_hd__mux2_2
XFILLER_0_86_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_952 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1222 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23130_ VGND VPWR VPWR VGND _02280_ _03509_ _03510_ _06976_ _07045_ sky130_fd_sc_hd__o31a_2
XFILLER_0_31_527 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20342_ VGND VPWR _00940_ _05597_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_82_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_909 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23061_ VPWR VGND VPWR VGND _06924_ _03293_ _03291_ _03794_ _03290_ _07004_ sky130_fd_sc_hd__a221o_2
X_20273_ VGND VPWR _00907_ _05561_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22012_ VPWR VGND keymem.key_mem\[3\]\[69\] _06487_ _06484_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_256_942 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_122_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_209_891 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_97_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23963_ VGND VPWR VPWR VGND clk _00456_ reset_n keymem.key_mem\[13\]\[84\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25702_ keymem.prev_key1_reg\[18\] clk _02195_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_93_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22914_ VGND VPWR _06914_ _06880_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_58_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23894_ VGND VPWR VPWR VGND clk _00387_ reset_n keymem.key_mem\[13\]\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25633_ VGND VPWR VPWR VGND clk _02126_ reset_n keymem.key_mem\[0\]\[90\] sky130_fd_sc_hd__dfrtp_2
X_22845_ VPWR VGND VPWR VGND keymem.rcon_logic.tmp_rcon\[6\] _06864_ keymem.rcon_logic.tmp_rcon\[7\]
+ _06867_ _02170_ sky130_fd_sc_hd__a22o_2
XFILLER_0_252_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25564_ VGND VPWR VPWR VGND clk _02057_ reset_n keymem.key_mem\[0\]\[21\] sky130_fd_sc_hd__dfrtp_2
X_22776_ VGND VPWR _06850_ _06779_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24515_ VGND VPWR VPWR VGND clk _01008_ reset_n keymem.key_mem\[9\]\[124\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_133_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21727_ VGND VPWR _01589_ _06333_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25495_ VGND VPWR VPWR VGND clk _01988_ reset_n keymem.key_mem\[1\]\[80\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_30_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24446_ VGND VPWR VPWR VGND clk _00939_ reset_n keymem.key_mem\[9\]\[55\] sky130_fd_sc_hd__dfrtp_2
X_12460_ VGND VPWR _08032_ _07685_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21658_ VGND VPWR _06297_ _06262_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_168_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_34_321 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_164_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20609_ VGND VPWR _01066_ _05738_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12391_ VGND VPWR _07969_ _07557_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24377_ VGND VPWR VPWR VGND clk _00870_ reset_n keymem.key_mem\[10\]\[114\] sky130_fd_sc_hd__dfrtp_2
X_21589_ VGND VPWR _01524_ _06260_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_151_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_65_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14130_ VGND VPWR _09600_ _09336_ _09601_ _09343_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_23328_ VPWR VGND VGND VPWR _07206_ _07207_ _04382_ sky130_fd_sc_hd__nor2_2
XFILLER_0_244_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_104_275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_240_1317 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14061_ VGND VPWR _09533_ _07378_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_244_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23259_ VPWR VGND VPWR VGND _07144_ block[5] _04837_ enc_block.block_w2_reg\[5\]
+ _04798_ _07145_ sky130_fd_sc_hd__a221o_2
X_13012_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[84\] _08449_ _08530_ _08526_ _08531_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_105_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17820_ VGND VPWR VPWR VGND _03777_ _03808_ keymem.prev_key0_reg\[66\] _03809_ sky130_fd_sc_hd__mux2_2
XFILLER_0_101_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_400 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_175_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17751_ VGND VPWR VPWR VGND _03763_ _02961_ keymem.prev_key0_reg\[41\] _03765_ sky130_fd_sc_hd__mux2_2
X_14963_ VGND VPWR VGND VPWR enc_block.block_w2_reg\[14\] _09269_ _09021_ _10425_
+ _10427_ _10426_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_55_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_175_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16702_ VGND VPWR VGND VPWR _02853_ keymem.prev_key1_reg\[95\] _02855_ _02852_ sky130_fd_sc_hd__nand3_2
X_13914_ VGND VPWR _09386_ _09318_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_215_861 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17682_ VGND VPWR VPWR VGND _03703_ _03717_ keymem.prev_key0_reg\[19\] _03718_ sky130_fd_sc_hd__mux2_2
X_14894_ VGND VPWR VGND VPWR _10349_ _10358_ _10359_ _10345_ _10357_ sky130_fd_sc_hd__nor4_2
XFILLER_0_18_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19421_ VPWR VGND keymem.key_mem\[12\]\[10\] _05107_ _05102_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16633_ VGND VPWR _00040_ _02788_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13845_ VGND VPWR _09317_ _09316_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_230_853 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_18_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_216_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_162_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_71_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19352_ VPWR VGND keymem.key_mem_we _05062_ _03580_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16564_ VGND VPWR _00037_ _02722_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_186_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_155_2_Right_227 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13776_ VGND VPWR _09248_ _09247_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18303_ VPWR VGND VGND VPWR _04204_ enc_block.block_w2_reg\[12\] enc_block.block_w2_reg\[13\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_112_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15515_ VGND VPWR VGND VPWR _10973_ _10974_ _10966_ _10964_ _10975_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_84_243 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12727_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[56\] _07748_ keymem.key_mem\[11\]\[56\]
+ _08090_ _08274_ sky130_fd_sc_hd__a22o_2
X_19283_ VPWR VGND keymem.key_mem\[13\]\[90\] _05017_ _04979_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16495_ VPWR VGND VGND VPWR _02655_ _02656_ _02654_ sky130_fd_sc_hd__nor2_2
X_18234_ VGND VPWR _04141_ enc_block.block_w3_reg\[7\] enc_block.block_w2_reg\[14\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15446_ VGND VPWR VGND VPWR _09523_ _10905_ _10903_ _10904_ _10907_ sky130_fd_sc_hd__a31o_2
X_12658_ VGND VPWR _08211_ _07903_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_37_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_53_630 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_182_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_343 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18165_ VGND VPWR _04078_ enc_block.block_w3_reg\[1\] _03985_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15377_ VGND VPWR _10838_ _08928_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_13_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12589_ VGND VPWR VGND VPWR _07584_ keymem.key_mem\[14\]\[43\] _08146_ _08148_ _08149_
+ _08069_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_154_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_105_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17116_ VGND VPWR VPWR VGND _03230_ _03231_ keymem.prev_key0_reg\[69\] _10189_ _10187_
+ sky130_fd_sc_hd__a31oi_2
XFILLER_0_20_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14328_ VPWR VGND VGND VPWR _09033_ _09798_ _09148_ sky130_fd_sc_hd__nor2_2
XFILLER_0_68_1183 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18096_ VPWR VGND VGND VPWR _04015_ _04010_ _04013_ sky130_fd_sc_hd__nand2_2
XFILLER_0_262_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_900 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_111_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_13 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_223_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17047_ VGND VPWR VGND VPWR _02832_ _02831_ _03169_ keymem.prev_key1_reg\[62\] sky130_fd_sc_hd__a21oi_2
XFILLER_0_29_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14259_ VGND VPWR _09729_ _08926_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_988 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_999 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_29_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_267_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_209_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18998_ VPWR VGND VGND VPWR _04778_ _04829_ _04248_ sky130_fd_sc_hd__nor2_2
XFILLER_0_178_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17949_ VGND VPWR _00247_ _03897_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_206_850 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_136_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20960_ VGND VPWR VPWR VGND _05912_ _05015_ keymem.key_mem\[7\]\[89\] _05927_ sky130_fd_sc_hd__mux2_2
XFILLER_0_139_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19619_ VGND VPWR _00602_ _05212_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_205_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20891_ VGND VPWR VGND VPWR _05890_ keymem.key_mem_we _03109_ _05864_ _01196_ sky130_fd_sc_hd__a31o_2
XFILLER_0_36_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22630_ VGND VPWR VPWR VGND _06785_ keymem.key_mem\[0\]\[4\] _10099_ _06786_ sky130_fd_sc_hd__mux2_2
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_105_2_Left_576 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22561_ VGND VPWR _01991_ _06765_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_265 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_61_82 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_1_Left_341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_75_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21512_ VGND VPWR VPWR VGND _06209_ _03443_ keymem.key_mem\[5\]\[93\] _06219_ sky130_fd_sc_hd__mux2_2
X_24300_ VGND VPWR VPWR VGND clk _00793_ reset_n keymem.key_mem\[10\]\[37\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_3_Right_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_118_356 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_267_1453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22492_ VGND VPWR _06737_ _06696_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_228_1404 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25280_ VGND VPWR VPWR VGND clk _01773_ reset_n keymem.key_mem\[3\]\[121\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_855 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_118_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_8_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21443_ VGND VPWR VPWR VGND _06173_ _03149_ keymem.key_mem\[5\]\[60\] _06183_ sky130_fd_sc_hd__mux2_2
X_24231_ VGND VPWR VPWR VGND clk _00724_ reset_n keymem.key_mem\[11\]\[96\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_267_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24162_ VGND VPWR VPWR VGND clk _00655_ reset_n keymem.key_mem\[11\]\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_847 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_86_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21374_ VGND VPWR VPWR VGND _06140_ _02764_ keymem.key_mem\[5\]\[27\] _06147_ sky130_fd_sc_hd__mux2_2
XFILLER_0_32_858 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_32_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23113_ VGND VPWR _02273_ _07035_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20325_ VGND VPWR _00932_ _05588_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24093_ VGND VPWR VPWR VGND clk _00586_ reset_n keymem.key_mem\[12\]\[86\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_261_1096 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23044_ VGND VPWR _02246_ _06993_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20256_ VGND VPWR _00899_ _05552_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20187_ VGND VPWR VPWR VGND _05504_ _03573_ keymem.key_mem\[10\]\[113\] _05514_ sky130_fd_sc_hd__mux2_2
XFILLER_0_157_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24995_ VGND VPWR VPWR VGND clk _01488_ reset_n keymem.key_mem\[5\]\[92\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_243_466 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_157_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23946_ VGND VPWR VPWR VGND clk _00439_ reset_n keymem.key_mem\[13\]\[67\] sky130_fd_sc_hd__dfrtp_2
X_11960_ VPWR VGND VGND VPWR _07548_ _07563_ _07543_ sky130_fd_sc_hd__nor2_2
XFILLER_0_118_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11891_ VGND VPWR result[112] _07509_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23877_ VGND VPWR VPWR VGND clk _00370_ reset_n enc_block.block_w2_reg\[30\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_211_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_402 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13630_ VGND VPWR _09102_ _09101_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25616_ VGND VPWR VPWR VGND clk _02109_ reset_n keymem.key_mem\[0\]\[73\] sky130_fd_sc_hd__dfrtp_2
X_22828_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[127\] _06839_ _03864_ _05089_ _02163_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_170_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13561_ VGND VPWR _09033_ _09032_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_109_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25547_ VGND VPWR VPWR VGND clk _02040_ reset_n keymem.key_mem\[0\]\[4\] sky130_fd_sc_hd__dfrtp_2
X_22759_ VPWR VGND VGND VPWR _06844_ keymem.key_mem\[0\]\[75\] _06839_ sky130_fd_sc_hd__nand2_2
X_15300_ VPWR VGND VGND VPWR _10538_ _10762_ _10628_ sky130_fd_sc_hd__nor2_2
X_12512_ VPWR VGND VPWR VGND _08078_ keymem.key_mem\[5\]\[36\] _07725_ keymem.key_mem\[4\]\[36\]
+ _08077_ _08079_ sky130_fd_sc_hd__a221o_2
X_16280_ VPWR VGND VPWR VGND _11410_ _11513_ _11435_ _11260_ _02444_ sky130_fd_sc_hd__or4_2
XFILLER_0_81_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13492_ VGND VPWR _08964_ _08941_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25478_ VGND VPWR VPWR VGND clk _01971_ reset_n keymem.key_mem\[1\]\[63\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_240_Right_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_212_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_168_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15231_ VPWR VGND VGND VPWR _10462_ _10467_ _10694_ _10521_ _10469_ sky130_fd_sc_hd__o22ai_2
X_12443_ VGND VPWR _08016_ _07609_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24429_ VGND VPWR VPWR VGND clk _00922_ reset_n keymem.key_mem\[9\]\[38\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_99_2_Left_570 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_129_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_136_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_836 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_65_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15162_ VPWR VGND VPWR VGND _10625_ _10626_ _10622_ _10624_ sky130_fd_sc_hd__or3b_2
XFILLER_0_22_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12374_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[24\] _07779_ keymem.key_mem\[3\]\[24\]
+ _07603_ _07953_ sky130_fd_sc_hd__a22o_2
X_14113_ VPWR VGND VPWR VGND _09580_ _09583_ _09581_ _09579_ _09584_ sky130_fd_sc_hd__or4_2
XFILLER_0_65_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1114 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15093_ VGND VPWR _10557_ _10556_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19970_ VGND VPWR _05400_ _05388_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_132_392 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_205_1245 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18921_ VPWR VGND _04760_ _04759_ enc_block.round_key\[49\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_14044_ VGND VPWR _09516_ _09515_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_157_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_24_1075 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18852_ VPWR VGND VPWR VGND _04697_ block[42] _04576_ enc_block.block_w0_reg\[10\]
+ _04666_ _04698_ sky130_fd_sc_hd__a221o_2
XFILLER_0_237_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17803_ VGND VPWR VGND VPWR _03732_ keymem.prev_key1_reg\[60\] _03798_ _03789_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_175_1311 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18783_ VPWR VGND _04635_ enc_block.block_w1_reg\[7\] enc_block.block_w1_reg\[3\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_15995_ VGND VPWR VGND VPWR _10728_ _10677_ _11450_ keymem.prev_key1_reg\[113\] sky130_fd_sc_hd__a21oi_2
XFILLER_0_179_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_915 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17734_ VGND VPWR VPWR VGND _03723_ _02887_ keymem.prev_key0_reg\[34\] _03755_ sky130_fd_sc_hd__mux2_2
X_14946_ VPWR VGND VPWR VGND _10397_ _10409_ _10403_ _10392_ _10410_ sky130_fd_sc_hd__or4_2
XFILLER_0_261_263 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_82_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_262_797 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_76_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17665_ VGND VPWR _00154_ _03706_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14877_ VGND VPWR VGND VPWR _08999_ _09019_ _09177_ _09090_ _10341_ _10342_ sky130_fd_sc_hd__o32a_2
XFILLER_0_82_59 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_203_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_89_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_352 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16616_ VGND VPWR _02772_ keymem.prev_key0_reg\[60\] keymem.prev_key0_reg\[92\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
X_19404_ VPWR VGND keymem.key_mem\[12\]\[2\] _05098_ _05095_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13828_ VGND VPWR _09300_ _09266_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17596_ VGND VPWR VPWR VGND _03593_ keymem.key_mem\[14\]\[125\] _03654_ _03655_ sky130_fd_sc_hd__mux2_2
XFILLER_0_203_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_202_374 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_230_694 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_212_1238 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_1171 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_159_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19335_ VGND VPWR VPWR VGND _05046_ _05050_ keymem.key_mem\[13\]\[108\] _05051_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_156_2_Right_228 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16547_ VPWR VGND VPWR VGND _02706_ key[25] _09719_ sky130_fd_sc_hd__or2_2
X_13759_ VGND VPWR VGND VPWR _09157_ _09029_ _09108_ _09156_ _09230_ _09231_ sky130_fd_sc_hd__o32a_2
XFILLER_0_174_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19266_ VPWR VGND keymem.key_mem_we _05006_ _03364_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16478_ VPWR VGND VPWR VGND _02639_ keymem.prev_key0_reg\[119\] sky130_fd_sc_hd__inv_2
XFILLER_0_122_54 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18217_ VGND VPWR VPWR VGND _03974_ enc_block.block_w0_reg\[13\] _04125_ _04126_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_186_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15429_ VGND VPWR VGND VPWR _10890_ _10482_ _10646_ _10667_ _10562_ sky130_fd_sc_hd__a211o_2
X_19197_ VPWR VGND keymem.key_mem\[13\]\[56\] _04965_ _04961_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_182_1304 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_147_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_348 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18148_ VPWR VGND VGND VPWR _04062_ _04063_ _04041_ sky130_fd_sc_hd__nor2_2
XFILLER_0_83_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18079_ VPWR VGND VGND VPWR _03999_ _03996_ _03998_ sky130_fd_sc_hd__nand2_2
XFILLER_0_44_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_514 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_40_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20110_ VGND VPWR VPWR VGND _05469_ _03295_ keymem.key_mem\[10\]\[76\] _05474_ sky130_fd_sc_hd__mux2_2
X_21090_ VGND VPWR VPWR VGND _05996_ _02549_ keymem.key_mem\[6\]\[21\] _05997_ sky130_fd_sc_hd__mux2_2
XFILLER_0_1_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_569 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20041_ VGND VPWR VPWR VGND _05435_ _02985_ keymem.key_mem\[10\]\[43\] _05438_ sky130_fd_sc_hd__mux2_2
XFILLER_0_42_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_265_580 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_147_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_158_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23800_ VGND VPWR VPWR VGND clk _00293_ reset_n enc_block.block_w0_reg\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24780_ VGND VPWR VPWR VGND clk _01273_ reset_n keymem.key_mem\[6\]\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_241_948 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21992_ VGND VPWR VGND VPWR _06476_ keymem.key_mem_we _03140_ _06475_ _01711_ sky130_fd_sc_hd__a31o_2
XFILLER_0_94_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23731_ keymem.prev_key0_reg\[87\] clk _00228_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20943_ VGND VPWR VGND VPWR _05918_ keymem.key_mem_we _03330_ _05916_ _01220_ sky130_fd_sc_hd__a31o_2
XFILLER_0_234_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_711 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_55_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23662_ keymem.prev_key0_reg\[18\] clk _00159_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_234_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20874_ VGND VPWR _01188_ _05881_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_163_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_49_755 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25401_ VGND VPWR VPWR VGND clk _01894_ reset_n keymem.key_mem\[2\]\[114\] sky130_fd_sc_hd__dfrtp_2
X_22613_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[123\] _06756_ _03793_ _05081_ _02031_
+ sky130_fd_sc_hd__a22o_2
X_23593_ VGND VPWR VPWR VGND clk _00094_ reset_n keymem.key_mem\[14\]\[82\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25332_ VGND VPWR VPWR VGND clk _01825_ reset_n keymem.key_mem\[2\]\[45\] sky130_fd_sc_hd__dfrtp_2
X_22544_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[72\] _06754_ _06753_ _04986_ _01980_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_64_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25263_ VGND VPWR VPWR VGND clk _01756_ reset_n keymem.key_mem\[3\]\[104\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_173_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_118_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22475_ VGND VPWR VPWR VGND _06726_ keymem.key_mem\[1\]\[31\] _02862_ _06732_ sky130_fd_sc_hd__mux2_2
XFILLER_0_165_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_359 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_133_134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24214_ VGND VPWR VPWR VGND clk _00707_ reset_n keymem.key_mem\[11\]\[79\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_133_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21426_ VGND VPWR _01447_ _06174_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_126_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25194_ VGND VPWR VPWR VGND clk _01687_ reset_n keymem.key_mem\[3\]\[35\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_71_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_206_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21357_ VGND VPWR VPWR VGND _06128_ _02409_ keymem.key_mem\[5\]\[19\] _06138_ sky130_fd_sc_hd__mux2_2
X_24145_ VGND VPWR VPWR VGND clk _00638_ reset_n keymem.key_mem\[11\]\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_241_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20308_ VGND VPWR _00924_ _05579_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_198_1311 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12090_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[4\] _07534_ _07688_ _07682_ _07689_
+ sky130_fd_sc_hd__o22a_2
X_24076_ VGND VPWR VPWR VGND clk _00569_ reset_n keymem.key_mem\[12\]\[69\] sky130_fd_sc_hd__dfrtp_2
X_21288_ VGND VPWR _01383_ _06100_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_202_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20239_ VGND VPWR _00891_ _05543_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23027_ VPWR VGND VGND VPWR _06983_ _03178_ _06976_ sky130_fd_sc_hd__nand2_2
XFILLER_0_60_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_239_1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14800_ VGND VPWR VGND VPWR _10265_ _10263_ _10266_ _10264_ sky130_fd_sc_hd__nand3_2
XFILLER_0_244_786 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_216_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15780_ VGND VPWR _11236_ _11235_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_204_628 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12992_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[82\] _08449_ _08512_ _08506_ _08513_
+ sky130_fd_sc_hd__o22a_2
X_24978_ VGND VPWR VPWR VGND clk _01471_ reset_n keymem.key_mem\[5\]\[75\] sky130_fd_sc_hd__dfrtp_2
X_14731_ VGND VPWR VGND VPWR _09157_ _09068_ _09072_ _09124_ _10197_ sky130_fd_sc_hd__o22a_2
XFILLER_0_203_138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23929_ VGND VPWR VPWR VGND clk _00422_ reset_n keymem.key_mem\[13\]\[50\] sky130_fd_sc_hd__dfrtp_2
X_11943_ VGND VPWR _07546_ _07545_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_197_830 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_19_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17450_ VPWR VGND VGND VPWR _03528_ _10817_ _10818_ sky130_fd_sc_hd__nand2_2
X_14662_ VPWR VGND VGND VPWR _09423_ _09330_ _09383_ _09355_ _10129_ _10128_ sky130_fd_sc_hd__o221a_2
XFILLER_0_52_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_210 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11874_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[8\] dec_new_block\[104\]
+ _07501_ sky130_fd_sc_hd__mux2_2
XFILLER_0_86_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16401_ VGND VPWR VGND VPWR _11493_ _11412_ _11224_ _11407_ _02563_ sky130_fd_sc_hd__a31o_2
XFILLER_0_200_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1480 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13613_ VPWR VGND VGND VPWR _09085_ _08958_ _09010_ sky130_fd_sc_hd__nand2_2
XFILLER_0_213_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17381_ VGND VPWR _00108_ _03468_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_156_226 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14593_ VPWR VGND VGND VPWR _09456_ _09358_ _10061_ _09350_ _09749_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_27_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19120_ VPWR VGND keymem.key_mem\[13\]\[28\] _04916_ _04915_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16332_ VGND VPWR VPWR VGND _02494_ _02483_ _02482_ _02495_ sky130_fd_sc_hd__mux2_2
X_13544_ VPWR VGND VPWR VGND _09014_ _09015_ _08991_ _08977_ _09016_ sky130_fd_sc_hd__or4_2
XFILLER_0_54_224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_109_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19051_ VPWR VGND VPWR VGND _04875_ _04874_ _04873_ enc_block.block_w2_reg\[31\]
+ _04613_ _00371_ sky130_fd_sc_hd__a221o_2
X_16263_ VPWR VGND VPWR VGND _11227_ _11460_ _11228_ _11226_ _02427_ sky130_fd_sc_hd__or4_2
XFILLER_0_42_408 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_2_Right_152 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13475_ VPWR VGND VPWR VGND _08947_ enc_block.sword_ctr_reg\[1\] sky130_fd_sc_hd__inv_2
X_18002_ VGND VPWR VGND VPWR _03737_ keymem.prev_key1_reg\[124\] _03933_ _03789_ sky130_fd_sc_hd__a21oi_2
X_15214_ VPWR VGND VGND VPWR _10493_ _10671_ _10676_ _10677_ sky130_fd_sc_hd__nor3_2
X_12426_ VGND VPWR VGND VPWR _08001_ _07908_ keymem.key_mem\[6\]\[28\] _07998_ _08000_
+ sky130_fd_sc_hd__a211o_2
X_16194_ VPWR VGND VGND VPWR _11372_ _02359_ _11464_ sky130_fd_sc_hd__nor2_2
XFILLER_0_22_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_50_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15145_ VGND VPWR _10609_ _10458_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12357_ VGND VPWR VGND VPWR _07838_ keymem.key_mem\[11\]\[22\] _07935_ _07937_ _07938_
+ _07662_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_26_1137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_267_834 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15076_ VPWR VGND VPWR VGND _10457_ _10435_ _10444_ _10419_ _10540_ sky130_fd_sc_hd__or4_2
XFILLER_0_77_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19953_ VGND VPWR _00757_ _05391_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12288_ VPWR VGND VPWR VGND _07873_ keymem.key_mem\[9\]\[17\] _07717_ keymem.key_mem\[11\]\[17\]
+ _07781_ _07874_ sky130_fd_sc_hd__a221o_2
X_14027_ VPWR VGND VGND VPWR _09293_ _09434_ _09499_ _09386_ _09443_ sky130_fd_sc_hd__o22ai_2
X_18904_ VGND VPWR _04744_ _03957_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_142_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_120_395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19884_ VGND VPWR _00726_ _05353_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18835_ VGND VPWR VGND VPWR _04681_ _04680_ _04682_ _00348_ sky130_fd_sc_hd__a21o_2
XFILLER_0_208_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18766_ _04618_ _04620_ _04560_ _04619_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_15978_ VGND VPWR VGND VPWR _11434_ _11273_ _11289_ _11227_ _11288_ sky130_fd_sc_hd__and4_2
XFILLER_0_93_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1152 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_26_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14929_ enc_block.sword_ctr_reg\[1\] _10393_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[8\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_17717_ VPWR VGND VPWR VGND _02762_ _03744_ keymem.prev_key0_reg\[27\] _03730_ _00168_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_37_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18697_ VPWR VGND _04558_ _04557_ enc_block.round_key\[91\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_26_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17648_ VGND VPWR VPWR VGND _03681_ _03694_ keymem.prev_key0_reg\[8\] _03695_ sky130_fd_sc_hd__mux2_2
XFILLER_0_212_1046 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17579_ VPWR VGND VPWR VGND _03639_ _03636_ _03635_ key[251] _08929_ _03640_ sky130_fd_sc_hd__a221o_2
XFILLER_0_46_725 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19318_ VPWR VGND keymem.key_mem_we _05039_ _03511_ VPWR VGND sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_157_2_Right_229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_85_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20590_ VGND VPWR _01057_ _05728_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_50_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19249_ VGND VPWR VPWR VGND _04993_ _04995_ keymem.key_mem\[13\]\[77\] _04996_ sky130_fd_sc_hd__mux2_2
XFILLER_0_5_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22260_ VGND VPWR _01837_ _06618_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_182_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_103_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21211_ VGND VPWR VPWR VGND _06052_ _03321_ keymem.key_mem\[6\]\[79\] _06060_ sky130_fd_sc_hd__mux2_2
XFILLER_0_258_801 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22191_ VGND VPWR _01804_ _06582_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_13_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_496 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21142_ VGND VPWR VPWR VGND _06018_ _03015_ keymem.key_mem\[6\]\[46\] _06024_ sky130_fd_sc_hd__mux2_2
XFILLER_0_160_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_160_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21073_ VGND VPWR VPWR VGND _05983_ _11039_ keymem.key_mem\[6\]\[13\] _05988_ sky130_fd_sc_hd__mux2_2
XFILLER_0_67_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20024_ VGND VPWR VPWR VGND _05424_ _02904_ keymem.key_mem\[10\]\[35\] _05429_ sky130_fd_sc_hd__mux2_2
X_24901_ VGND VPWR VPWR VGND clk _01394_ reset_n keymem.key_mem\[6\]\[126\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_253_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24832_ VGND VPWR VPWR VGND clk _01325_ reset_n keymem.key_mem\[6\]\[57\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24763_ VGND VPWR VPWR VGND clk _01256_ reset_n keymem.key_mem\[7\]\[116\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21975_ VGND VPWR VPWR VGND _06462_ _04958_ keymem.key_mem\[3\]\[52\] _06467_ sky130_fd_sc_hd__mux2_2
XFILLER_0_174_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_197_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23714_ keymem.prev_key0_reg\[70\] clk _00211_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20926_ VPWR VGND keymem.key_mem\[7\]\[73\] _05909_ _05899_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_178_351 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24694_ VGND VPWR VPWR VGND clk _01187_ reset_n keymem.key_mem\[7\]\[47\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_95_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_178_384 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23645_ keymem.prev_key0_reg\[1\] clk _00142_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20857_ VGND VPWR _01180_ _05872_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_260_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23576_ VGND VPWR VPWR VGND clk _00077_ reset_n keymem.key_mem\[14\]\[65\] sky130_fd_sc_hd__dfrtp_2
X_20788_ VPWR VGND keymem.key_mem\[7\]\[9\] _05835_ _05830_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_14_1085 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25315_ VGND VPWR VPWR VGND clk _01808_ reset_n keymem.key_mem\[2\]\[28\] sky130_fd_sc_hd__dfrtp_2
X_22527_ VGND VPWR _01971_ _06751_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25246_ VGND VPWR VPWR VGND clk _01739_ reset_n keymem.key_mem\[3\]\[87\] sky130_fd_sc_hd__dfrtp_2
X_13260_ VPWR VGND VPWR VGND _08753_ keymem.key_mem\[9\]\[109\] _07672_ keymem.key_mem\[10\]\[109\]
+ _07876_ _08754_ sky130_fd_sc_hd__a221o_2
X_22458_ VGND VPWR VPWR VGND _06715_ keymem.key_mem\[1\]\[23\] _02661_ _06723_ sky130_fd_sc_hd__mux2_2
XFILLER_0_33_953 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_106_178 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_66_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_27_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_975 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12211_ VPWR VGND VPWR VGND _07802_ keymem.key_mem\[13\]\[11\] _07587_ keymem.key_mem\[11\]\[11\]
+ _07761_ _07803_ sky130_fd_sc_hd__a221o_2
X_21409_ VGND VPWR _01439_ _06165_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13191_ VPWR VGND VPWR VGND _08691_ keymem.key_mem\[9\]\[102\] _07716_ keymem.key_mem\[10\]\[102\]
+ _08193_ _08692_ sky130_fd_sc_hd__a221o_2
X_25177_ VGND VPWR VPWR VGND clk _01670_ reset_n keymem.key_mem\[3\]\[18\] sky130_fd_sc_hd__dfrtp_2
X_22389_ VGND VPWR VPWR VGND _06680_ _03613_ keymem.key_mem\[2\]\[119\] _06686_ sky130_fd_sc_hd__mux2_2
XFILLER_0_27_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12142_ VGND VPWR _07738_ _07591_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24128_ VGND VPWR VPWR VGND clk _00621_ reset_n keymem.key_mem\[12\]\[121\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_206_1373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_21_1001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16950_ VGND VPWR VGND VPWR _03079_ _03080_ _03078_ keylen _03081_ sky130_fd_sc_hd__a2bb2o_2
X_24059_ VGND VPWR VPWR VGND clk _00552_ reset_n keymem.key_mem\[12\]\[52\] sky130_fd_sc_hd__dfrtp_2
X_12073_ VGND VPWR _07673_ _07577_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_25_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15901_ VGND VPWR VGND VPWR _11357_ _11208_ _11228_ _11272_ _11288_ sky130_fd_sc_hd__and4_2
XFILLER_0_21_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16881_ VGND VPWR VPWR VGND _10091_ key[175] keymem.prev_key1_reg\[47\] _03018_ sky130_fd_sc_hd__mux2_2
XFILLER_0_232_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_159_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15832_ VGND VPWR _11288_ _11187_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18620_ VGND VPWR _04489_ enc_block.block_w2_reg\[23\] enc_block.block_w1_reg\[27\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_745 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15763_ VGND VPWR _11219_ _11218_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18551_ VPWR VGND _04427_ enc_block.block_w3_reg\[15\] enc_block.block_w3_reg\[11\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_63_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12975_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[81\] _07812_ keymem.key_mem\[10\]\[81\]
+ _08193_ _08497_ sky130_fd_sc_hd__a22o_2
XFILLER_0_204_469 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_38_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_789 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14714_ VGND VPWR VGND VPWR _09020_ _09105_ _10179_ _09938_ _10181_ _10180_ sky130_fd_sc_hd__a2111o_2
X_17502_ VGND VPWR VGND VPWR _03152_ key[241] _03572_ _03573_ sky130_fd_sc_hd__a21o_2
XFILLER_0_86_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18482_ VGND VPWR _04365_ enc_block.block_w0_reg\[4\] _04364_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_11926_ VGND VPWR VPWR VGND encdec enc_block.round\[2\] dec_round_nr\[2\] _07529_
+ sky130_fd_sc_hd__mux2_2
X_15694_ VGND VPWR _00027_ _11150_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17433_ VGND VPWR VPWR VGND _03029_ _10655_ key[104] _03513_ sky130_fd_sc_hd__mux2_2
X_14645_ VPWR VGND VPWR VGND _09499_ _10111_ _10112_ _09482_ _09496_ sky130_fd_sc_hd__or4b_2
X_11857_ VGND VPWR result[95] _07492_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_67_371 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17364_ VGND VPWR _00106_ _03453_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_248_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14576_ VGND VPWR VGND VPWR _09476_ _09399_ _09576_ _10044_ sky130_fd_sc_hd__a21o_2
X_11788_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[29\] dec_new_block\[61\]
+ _07458_ sky130_fd_sc_hd__mux2_2
XFILLER_0_248_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16315_ VPWR VGND VPWR VGND _02478_ _10085_ _02468_ key[148] _11043_ _02479_ sky130_fd_sc_hd__a221o_2
X_19103_ VGND VPWR VGND VPWR _04906_ keymem.key_mem_we _02480_ _04896_ _00392_ sky130_fd_sc_hd__a31o_2
X_13527_ VGND VPWR _08999_ _08998_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17295_ VGND VPWR VGND VPWR _03392_ _03152_ key[215] _03387_ _03391_ sky130_fd_sc_hd__a211o_2
XFILLER_0_137_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19034_ VGND VPWR _04860_ _04283_ _00369_ _04602_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_36_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_2_Right_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_109_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16246_ VGND VPWR VPWR VGND _11041_ keymem.key_mem\[14\]\[19\] _02410_ _02411_ sky130_fd_sc_hd__mux2_2
X_13458_ VGND VPWR _08930_ _08929_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_148_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_964 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12409_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[27\] _07596_ keymem.key_mem\[1\]\[27\]
+ _07557_ _07985_ sky130_fd_sc_hd__a22o_2
X_16177_ VGND VPWR _02342_ _09795_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13389_ VGND VPWR VGND VPWR _07841_ keymem.key_mem\[4\]\[122\] _08867_ _08869_ _08870_
+ _07573_ sky130_fd_sc_hd__a2111o_2
X_15128_ VPWR VGND VPWR VGND _10473_ _10409_ _10452_ _10439_ _10592_ sky130_fd_sc_hd__or4_2
XFILLER_0_259_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15059_ VPWR VGND VGND VPWR _10496_ _10519_ _10523_ _10522_ _10520_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_255_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_259_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19936_ VGND VPWR _00751_ _05380_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_114_2_Left_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_103_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19867_ VGND VPWR _00718_ _05344_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_37_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_83_1_Left_350 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_235_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18818_ VGND VPWR _04667_ enc_block.block_w2_reg\[30\] enc_block.block_w0_reg\[15\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_253_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19798_ VGND VPWR _00685_ _05308_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_74_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_194_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_211_907 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18749_ VGND VPWR _04604_ enc_block.block_w2_reg\[31\] enc_block.block_w0_reg\[9\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_204_970 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_144_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_204_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21760_ VGND VPWR _01605_ _06350_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_144_74 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20711_ VGND VPWR _01115_ _05791_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_187_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_153_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_714 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_92_105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21691_ VGND VPWR _01572_ _06314_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_50_1230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23430_ VPWR VGND VGND VPWR _07298_ enc_block.block_w3_reg\[31\] enc_block.block_w1_reg\[14\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_46_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20642_ VGND VPWR _01082_ _05755_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_11_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23361_ VPWR VGND _07237_ _07236_ enc_block.round_key\[15\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_20573_ VGND VPWR _01049_ _05719_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_2_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25100_ VGND VPWR VPWR VGND clk _01593_ reset_n keymem.key_mem\[4\]\[69\] sky130_fd_sc_hd__dfrtp_2
X_22312_ VGND VPWR _01862_ _06645_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_6_674 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23292_ VGND VPWR VGND VPWR _07173_ _03992_ _07174_ _02313_ sky130_fd_sc_hd__a21o_2
XFILLER_0_85_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_264_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_249_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25031_ VGND VPWR VPWR VGND clk _01524_ reset_n keymem.key_mem\[4\]\[0\] sky130_fd_sc_hd__dfrtp_2
X_22243_ VGND VPWR _01829_ _06609_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22174_ VGND VPWR _01796_ _06573_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_203_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_826 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_257_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21125_ VGND VPWR VPWR VGND _06007_ _02934_ keymem.key_mem\[6\]\[38\] _06015_ sky130_fd_sc_hd__mux2_2
XFILLER_0_121_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_160_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21056_ VGND VPWR _01273_ _05978_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_121_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20007_ VGND VPWR VPWR VGND _05413_ _02765_ keymem.key_mem\[10\]\[27\] _05420_ sky130_fd_sc_hd__mux2_2
XFILLER_0_214_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_92_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24815_ VGND VPWR VPWR VGND clk _01308_ reset_n keymem.key_mem\[6\]\[40\] sky130_fd_sc_hd__dfrtp_2
X_25795_ keymem.prev_key1_reg\[111\] clk _02288_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_119_1186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12760_ VGND VPWR VGND VPWR _07588_ keymem.key_mem\[13\]\[59\] _08301_ _08303_ _08304_
+ _07573_ sky130_fd_sc_hd__a2111o_2
X_24746_ VGND VPWR VPWR VGND clk _01239_ reset_n keymem.key_mem\[7\]\[99\] sky130_fd_sc_hd__dfrtp_2
X_21958_ VGND VPWR VPWR VGND _06449_ _04943_ keymem.key_mem\[3\]\[44\] _06458_ sky130_fd_sc_hd__mux2_2
X_11711_ VGND VPWR result[22] _07419_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_132_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20909_ VGND VPWR VGND VPWR _05900_ keymem.key_mem_we _03194_ _05893_ _01204_ sky130_fd_sc_hd__a31o_2
XFILLER_0_171_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12691_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[53\] _07843_ keymem.key_mem\[6\]\[53\]
+ _07639_ _08241_ sky130_fd_sc_hd__a22o_2
X_24677_ VGND VPWR VPWR VGND clk _01170_ reset_n keymem.key_mem\[7\]\[30\] sky130_fd_sc_hd__dfrtp_2
X_21889_ VPWR VGND keymem.key_mem\[3\]\[12\] _06421_ _06413_ VPWR VGND sky130_fd_sc_hd__and2_2
X_14430_ VGND VPWR VGND VPWR _09899_ _09897_ _09749_ _09355_ _09898_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_132_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11642_ VPWR VGND VGND VPWR _07381_ enc_block.enc_ctrl_reg\[3\] _07380_ sky130_fd_sc_hd__nand2_2
X_23628_ VGND VPWR VPWR VGND clk _00129_ reset_n keymem.key_mem\[14\]\[117\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_166_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14361_ VPWR VGND VPWR VGND _09829_ _09830_ _09831_ _09180_ _09828_ sky130_fd_sc_hd__or4b_2
X_23559_ VGND VPWR VPWR VGND clk _00060_ reset_n keymem.key_mem\[14\]\[48\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_52_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16100_ VGND VPWR VGND VPWR _10814_ keymem.prev_key1_reg\[114\] _11554_ _10775_ sky130_fd_sc_hd__nand3_2
XFILLER_0_134_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13312_ VPWR VGND VPWR VGND _08800_ keymem.key_mem\[13\]\[114\] _08125_ keymem.key_mem\[1\]\[114\]
+ _07671_ _08801_ sky130_fd_sc_hd__a221o_2
XFILLER_0_24_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17080_ VGND VPWR VGND VPWR _03199_ _02928_ _02927_ key[65] sky130_fd_sc_hd__o21a_2
X_14292_ VPWR VGND VGND VPWR _09348_ _09357_ _09762_ _09294_ _09378_ sky130_fd_sc_hd__o22ai_2
X_16031_ VPWR VGND VGND VPWR _11336_ _11486_ _11422_ sky130_fd_sc_hd__nor2_2
XFILLER_0_33_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25229_ VGND VPWR VPWR VGND clk _01722_ reset_n keymem.key_mem\[3\]\[70\] sky130_fd_sc_hd__dfrtp_2
X_13243_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[107\] _08391_ keymem.key_mem\[8\]\[107\]
+ _07903_ _08739_ sky130_fd_sc_hd__a22o_2
XFILLER_0_126_1157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13174_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[100\] _08124_ _08676_ _08670_ _08677_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_143_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12125_ VGND VPWR _07722_ _07578_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_20_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17982_ VGND VPWR VPWR VGND _03674_ _03919_ keymem.prev_key0_reg\[117\] _03920_ sky130_fd_sc_hd__mux2_2
XFILLER_0_40_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_264_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_100_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19721_ VGND VPWR VPWR VGND _05259_ keymem.key_mem\[11\]\[21\] _02550_ _05268_ sky130_fd_sc_hd__mux2_2
X_16933_ VGND VPWR VGND VPWR _03063_ _03065_ _03061_ _03066_ _03058_ sky130_fd_sc_hd__o2bb2a_2
X_12056_ VGND VPWR _07656_ _07564_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_40_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_217_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_254_1400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19652_ VGND VPWR VPWR VGND _05227_ _05071_ keymem.key_mem\[12\]\[118\] _05230_ sky130_fd_sc_hd__mux2_2
X_16864_ VGND VPWR VPWR VGND _09521_ key[173] keymem.prev_key1_reg\[45\] _03003_ sky130_fd_sc_hd__mux2_2
XFILLER_0_204_222 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18603_ VGND VPWR VGND VPWR _04474_ _04473_ _04472_ _04470_ sky130_fd_sc_hd__o21a_2
XFILLER_0_245_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15815_ VPWR VGND VGND VPWR _11270_ _11271_ _11262_ sky130_fd_sc_hd__nor2_2
XFILLER_0_260_862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19583_ VGND VPWR VPWR VGND _05183_ _05008_ keymem.key_mem\[12\]\[85\] _05194_ sky130_fd_sc_hd__mux2_2
X_16795_ VGND VPWR _10378_ keymem.prev_key1_reg\[39\] _02940_ keymem.prev_key1_reg\[71\]
+ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_245_73 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15746_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[21\] _10402_ _11202_ _09255_ _11200_
+ _11201_ sky130_fd_sc_hd__a32oi_2
X_18534_ VPWR VGND VGND VPWR _04411_ _04412_ _04077_ sky130_fd_sc_hd__nor2_2
XFILLER_0_99_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12958_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[79\] _07562_ keymem.key_mem\[8\]\[79\]
+ _07878_ _08482_ sky130_fd_sc_hd__a22o_2
X_11909_ VGND VPWR result[121] _07518_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_150_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15677_ VGND VPWR VGND VPWR _11134_ _11133_ _11132_ _11131_ _11130_ sky130_fd_sc_hd__and4_2
X_18465_ VGND VPWR VGND VPWR _04349_ _04266_ _04316_ _04350_ enc_block.block_w1_reg\[3\]
+ sky130_fd_sc_hd__o2bb2a_2
X_12889_ VGND VPWR VGND VPWR _08420_ _08150_ keymem.key_mem\[3\]\[72\] _08417_ _08419_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_111_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17416_ VGND VPWR VGND VPWR _03499_ _03496_ _03495_ _02919_ _03498_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_135_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_150_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14628_ VGND VPWR _10096_ _07378_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_51_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18396_ _04286_ _04288_ _04008_ _04287_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_28_544 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_114_88 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_111_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17347_ VGND VPWR VGND VPWR _03438_ _09637_ _10323_ key[221] sky130_fd_sc_hd__o21a_2
X_14559_ VGND VPWR VGND VPWR _10020_ _10019_ _10022_ _10026_ _10027_ _09951_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_3_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17278_ VGND VPWR VPWR VGND _02588_ _02589_ keymem.prev_key0_reg\[86\] _03376_ sky130_fd_sc_hd__or3_2
XFILLER_0_3_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_109_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_622 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19017_ VPWR VGND VPWR VGND _04845_ _04788_ _04844_ enc_block.block_w2_reg\[27\]
+ _04613_ _00367_ sky130_fd_sc_hd__a221o_2
X_16229_ VPWR VGND _02372_ _02394_ _02393_ VPWR VGND sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_82_2_Right_154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_261_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_772 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_70_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_666 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_227_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19919_ VGND VPWR _00743_ _05371_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_254_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22930_ VGND VPWR _06924_ _06883_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_97_208 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22861_ VGND VPWR _02177_ _06879_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_250_350 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24600_ VGND VPWR VPWR VGND clk _01093_ reset_n keymem.key_mem\[8\]\[81\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21812_ VGND VPWR VPWR VGND _06377_ _03533_ keymem.key_mem\[4\]\[106\] _06378_ sky130_fd_sc_hd__mux2_2
XFILLER_0_250_383 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25580_ VGND VPWR VPWR VGND clk _02073_ reset_n keymem.key_mem\[0\]\[37\] sky130_fd_sc_hd__dfrtp_2
X_22792_ VGND VPWR _02131_ _06856_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_39_809 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24531_ VGND VPWR VPWR VGND clk _01024_ reset_n keymem.key_mem\[8\]\[12\] sky130_fd_sc_hd__dfrtp_2
X_21743_ VGND VPWR _01597_ _06341_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_171_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_148_354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24462_ VGND VPWR VPWR VGND clk _00955_ reset_n keymem.key_mem\[9\]\[71\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_65_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1304 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21674_ VGND VPWR _01564_ _06305_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23413_ VGND VPWR _07283_ enc_block.block_w2_reg\[5\] enc_block.block_w0_reg\[20\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_503 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20625_ VGND VPWR _01074_ _05746_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24393_ VGND VPWR VPWR VGND clk _00886_ reset_n keymem.key_mem\[9\]\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_62_834 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23344_ VGND VPWR _02318_ _07221_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_73_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20556_ VGND VPWR _01041_ _05710_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23275_ VGND VPWR _07159_ enc_block.block_w3_reg\[30\] _07158_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20487_ VGND VPWR VPWR VGND _05534_ _03661_ keymem.key_mem\[9\]\[126\] _05673_ sky130_fd_sc_hd__mux2_2
XFILLER_0_28_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25014_ VGND VPWR VPWR VGND clk _01507_ reset_n keymem.key_mem\[5\]\[111\] sky130_fd_sc_hd__dfrtp_2
X_22226_ VGND VPWR VPWR VGND _06600_ _02964_ keymem.key_mem\[2\]\[41\] _06601_ sky130_fd_sc_hd__mux2_2
XFILLER_0_203_1310 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_259_984 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22157_ VGND VPWR VPWR VGND _06554_ _10746_ keymem.key_mem\[2\]\[9\] _06564_ sky130_fd_sc_hd__mux2_2
XFILLER_0_218_336 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21108_ VGND VPWR VPWR VGND _05996_ _02838_ keymem.key_mem\[6\]\[30\] _06006_ sky130_fd_sc_hd__mux2_2
X_22088_ VGND VPWR _01757_ _06526_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_22_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13930_ VPWR VGND VPWR VGND _09261_ _09245_ _09300_ _09297_ _09402_ sky130_fd_sc_hd__or4_2
XFILLER_0_261_637 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21039_ VGND VPWR VPWR VGND _05819_ _05089_ keymem.key_mem\[7\]\[127\] _05968_ sky130_fd_sc_hd__mux2_2
XFILLER_0_96_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1199 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13861_ VGND VPWR _09333_ _09332_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_9_1001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15600_ VPWR VGND VPWR VGND _10787_ _10560_ _11058_ _10717_ _10716_ sky130_fd_sc_hd__or4b_2
XFILLER_0_57_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12812_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[65\] _07902_ keymem.key_mem\[10\]\[65\]
+ _07785_ _08350_ sky130_fd_sc_hd__a22o_2
XFILLER_0_214_597 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16580_ _02736_ _02738_ _02735_ _02737_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_9_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13792_ VGND VPWR VGND VPWR enc_block.block_w1_reg\[25\] _08948_ _09022_ _09262_
+ _09264_ _09263_ sky130_fd_sc_hd__a2111o_2
X_25778_ keymem.prev_key1_reg\[94\] clk _02271_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_15531_ VGND VPWR VGND VPWR _10530_ _10545_ _10497_ _10587_ _10990_ sky130_fd_sc_hd__o22a_2
X_12743_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[58\] _07690_ keymem.key_mem\[7\]\[58\]
+ _07650_ _08288_ sky130_fd_sc_hd__a22o_2
X_24729_ VGND VPWR VPWR VGND clk _01222_ reset_n keymem.key_mem\[7\]\[82\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18250_ _04154_ _04156_ _04008_ _04155_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_15462_ VPWR VGND VPWR VGND _10885_ _10722_ _10721_ _10921_ _10922_ sky130_fd_sc_hd__or4_2
XFILLER_0_60_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12674_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[51\] _07984_ keymem.key_mem\[2\]\[51\]
+ _07816_ _08226_ sky130_fd_sc_hd__a22o_2
XFILLER_0_49_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17201_ VGND VPWR _00089_ _03307_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14413_ VGND VPWR VPWR VGND _09462_ _09881_ _09457_ _09882_ sky130_fd_sc_hd__or3_2
X_18181_ VPWR VGND VPWR VGND _04092_ block[106] _04076_ enc_block.block_w2_reg\[10\]
+ _04007_ _04093_ sky130_fd_sc_hd__a221o_2
X_11625_ VPWR VGND VPWR VGND _07366_ init sky130_fd_sc_hd__inv_2
XFILLER_0_5_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15393_ VPWR VGND VPWR VGND _10782_ _10853_ _10854_ _10567_ _10852_ sky130_fd_sc_hd__or4b_2
XFILLER_0_64_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17132_ VGND VPWR VPWR VGND _03185_ keymem.key_mem\[14\]\[70\] _03245_ _03246_ sky130_fd_sc_hd__mux2_2
X_14344_ VPWR VGND VGND VPWR _09174_ _09122_ _09814_ _09128_ _09053_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_128_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_1565 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_167_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_878 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_107_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_107_284 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_69_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17063_ VGND VPWR _03184_ _03183_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14275_ VGND VPWR VPWR VGND _09358_ _09336_ _09745_ _09744_ _09742_ sky130_fd_sc_hd__o211a_2
X_16014_ VGND VPWR _11469_ _11370_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13226_ VGND VPWR enc_block.round_key\[105\] _08723_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_100_46 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13157_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[99\] _07631_ keymem.key_mem\[2\]\[99\]
+ _07697_ _08661_ sky130_fd_sc_hd__a22o_2
XFILLER_0_0_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_249_494 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12108_ VGND VPWR _07706_ _07583_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_237_656 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_236_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_209_358 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17965_ VGND VPWR VGND VPWR _03564_ keymem.prev_key1_reg\[112\] _03908_ _10371_ sky130_fd_sc_hd__a21bo_2
X_13088_ VGND VPWR _08599_ _07746_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_40_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19704_ VGND VPWR _05259_ _05246_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_18_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16916_ VGND VPWR VGND VPWR _03049_ _09796_ _11560_ _11622_ _03050_ sky130_fd_sc_hd__a31o_2
X_12039_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[2\] _07639_ keymem.key_mem\[1\]\[2\]
+ _07624_ _07640_ sky130_fd_sc_hd__a22o_2
XFILLER_0_75_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_205_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17896_ VGND VPWR VGND VPWR _03736_ keymem.prev_key0_reg\[89\] _03861_ _03407_ _00230_
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_139_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19635_ VGND VPWR VPWR VGND _05216_ _05054_ keymem.key_mem\[12\]\[110\] _05221_ sky130_fd_sc_hd__mux2_2
X_16847_ VGND VPWR _00055_ _02987_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_75_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_252_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19566_ VGND VPWR VPWR VGND _05183_ _04995_ keymem.key_mem\[12\]\[77\] _05185_ sky130_fd_sc_hd__mux2_2
X_16778_ VGND VPWR VPWR VGND _02884_ keymem.key_mem\[14\]\[37\] _02924_ _02925_ sky130_fd_sc_hd__mux2_2
XFILLER_0_34_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18517_ VPWR VGND VPWR VGND _04396_ block[72] _04351_ enc_block.block_w3_reg\[8\]
+ _03954_ _04397_ sky130_fd_sc_hd__a221o_2
X_15729_ VGND VPWR VGND VPWR enc_block.block_w2_reg\[23\] _09269_ _10387_ _11183_
+ _11185_ _11184_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_47_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19497_ VGND VPWR VPWR VGND _05138_ _04945_ keymem.key_mem\[12\]\[45\] _05148_ sky130_fd_sc_hd__mux2_2
XFILLER_0_34_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18448_ VPWR VGND VPWR VGND _04334_ _04331_ _04333_ sky130_fd_sc_hd__or2_2
XFILLER_0_111_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_150_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_111_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18379_ VPWR VGND _04273_ _04272_ enc_block.round_key\[124\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_172_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20410_ VGND VPWR VPWR VGND _05627_ _03409_ keymem.key_mem\[9\]\[89\] _05633_ sky130_fd_sc_hd__mux2_2
XFILLER_0_86_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21390_ VGND VPWR _01430_ _06155_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_146_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20341_ VGND VPWR VPWR VGND _05591_ _03109_ keymem.key_mem\[9\]\[56\] _05597_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_964 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_2_Right_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23060_ VGND VPWR _02252_ _07003_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20272_ VGND VPWR VPWR VGND _05558_ _02661_ keymem.key_mem\[9\]\[23\] _05561_ sky130_fd_sc_hd__mux2_2
XFILLER_0_261_1289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22011_ VGND VPWR VPWR VGND _01720_ _06406_ _03226_ _08922_ _06486_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_59_82 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_109_1_Left_376 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23962_ VGND VPWR VPWR VGND clk _00455_ reset_n keymem.key_mem\[13\]\[83\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25701_ keymem.prev_key1_reg\[17\] clk _02194_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_97_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_192_1339 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22913_ VGND VPWR VGND VPWR _02401_ _02343_ _02408_ _06913_ sky130_fd_sc_hd__a21o_2
XFILLER_0_157_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Left_284 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_230_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23893_ VGND VPWR VPWR VGND clk _00386_ reset_n keymem.key_mem\[13\]\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_895 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25632_ VGND VPWR VPWR VGND clk _02125_ reset_n keymem.key_mem\[0\]\[89\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22844_ VPWR VGND VPWR VGND keymem.rcon_logic.tmp_rcon\[5\] _06864_ keymem.rcon_logic.tmp_rcon\[6\]
+ _06867_ _02169_ sky130_fd_sc_hd__a22o_2
XFILLER_0_116_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25563_ VGND VPWR VPWR VGND clk _02056_ reset_n keymem.key_mem\[0\]\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22775_ VGND VPWR _06849_ _03733_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24514_ VGND VPWR VPWR VGND clk _01007_ reset_n keymem.key_mem\[9\]\[123\] sky130_fd_sc_hd__dfrtp_2
X_21726_ VGND VPWR VPWR VGND _06330_ _03202_ keymem.key_mem\[4\]\[65\] _06333_ sky130_fd_sc_hd__mux2_2
X_25494_ VGND VPWR VPWR VGND clk _01987_ reset_n keymem.key_mem\[1\]\[79\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_148_184 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_139_2_Left_610 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24445_ VGND VPWR VPWR VGND clk _00938_ reset_n keymem.key_mem\[9\]\[54\] sky130_fd_sc_hd__dfrtp_2
X_21657_ VGND VPWR _01556_ _06296_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_30_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_46_171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_168_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_46_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20608_ VGND VPWR VPWR VGND _05736_ _03090_ keymem.key_mem\[8\]\[54\] _05738_ sky130_fd_sc_hd__mux2_2
X_12390_ VGND VPWR _07968_ _07593_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24376_ VGND VPWR VPWR VGND clk _00869_ reset_n keymem.key_mem\[10\]\[113\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_164_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21588_ VGND VPWR VPWR VGND _06259_ _09536_ keymem.key_mem\[4\]\[0\] _06260_ sky130_fd_sc_hd__mux2_2
X_23327_ VGND VPWR _07206_ _07203_ _07205_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20539_ VGND VPWR _01033_ _05701_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_244_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14060_ VGND VPWR VPWR VGND _09531_ _09525_ _09520_ _09532_ sky130_fd_sc_hd__mux2_2
X_23258_ VPWR VGND VGND VPWR _07143_ _07144_ _04382_ sky130_fd_sc_hd__nor2_2
X_13011_ VGND VPWR VGND VPWR _08530_ _07665_ keymem.key_mem\[4\]\[84\] _08527_ _08529_
+ sky130_fd_sc_hd__a211o_2
X_22209_ VGND VPWR VPWR VGND _06589_ _02883_ keymem.key_mem\[2\]\[33\] _06592_ sky130_fd_sc_hd__mux2_2
X_23189_ VGND VPWR VGND VPWR _03657_ _03656_ _03660_ _07082_ sky130_fd_sc_hd__a21o_2
XFILLER_0_197_1228 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_101_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_486 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14962_ VGND VPWR VGND VPWR _10426_ enc_block.sword_ctr_reg\[0\] enc_block.block_w1_reg\[14\]
+ enc_block.sword_ctr_reg\[1\] sky130_fd_sc_hd__and3b_2
XFILLER_0_175_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17750_ VGND VPWR _00181_ _03764_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_234_648 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_175_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16701_ VGND VPWR VGND VPWR _02853_ _02852_ keymem.prev_key1_reg\[95\] _02854_ sky130_fd_sc_hd__a21o_2
X_13913_ VGND VPWR VGND VPWR _09385_ _09376_ _09372_ _09341_ _09384_ sky130_fd_sc_hd__o211ai_2
X_14893_ VGND VPWR VGND VPWR _10358_ _09969_ _09181_ _09970_ _10160_ sky130_fd_sc_hd__a211o_2
X_17681_ VGND VPWR VPWR VGND _03691_ key[147] keymem.prev_key1_reg\[19\] _03717_ sky130_fd_sc_hd__mux2_2
XFILLER_0_255_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_1044 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19420_ VGND VPWR VGND VPWR _05106_ keymem.key_mem_we _10747_ _05093_ _00509_ sky130_fd_sc_hd__a31o_2
XFILLER_0_18_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13844_ VGND VPWR VGND VPWR _09316_ _09244_ _09243_ keymem.prev_key1_reg\[24\] _09003_
+ _09002_ sky130_fd_sc_hd__a32o_2
XFILLER_0_251_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16632_ VGND VPWR VPWR VGND _02662_ keymem.key_mem\[14\]\[28\] _02787_ _02788_ sky130_fd_sc_hd__mux2_2
XFILLER_0_134_1223 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_214_394 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_230_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_251_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19351_ VGND VPWR _00485_ _05061_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13775_ VGND VPWR _09247_ _09246_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_29_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16563_ VGND VPWR VPWR VGND _02662_ keymem.key_mem\[14\]\[25\] _02721_ _02722_ sky130_fd_sc_hd__mux2_2
XFILLER_0_186_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18302_ VPWR VGND _04203_ _04045_ enc_block.block_w1_reg\[20\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_242_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12726_ VGND VPWR VGND VPWR _07908_ keymem.key_mem\[6\]\[56\] _08270_ _08272_ _08273_
+ _08243_ sky130_fd_sc_hd__a2111o_2
X_15514_ VGND VPWR VPWR VGND _10974_ _10278_ _10970_ _10969_ _07378_ sky130_fd_sc_hd__o31a_2
X_16494_ VGND VPWR VGND VPWR _09521_ _02653_ _02651_ _02652_ _02655_ sky130_fd_sc_hd__a31o_2
X_19282_ VGND VPWR _00461_ _05016_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_112_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18233_ VPWR VGND _04140_ enc_block.block_w0_reg\[31\] enc_block.block_w1_reg\[23\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_15445_ VGND VPWR VGND VPWR _10904_ _10903_ _10906_ _10905_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_123_2_Left_594 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12657_ VGND VPWR enc_block.round_key\[49\] _08210_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_37_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_706 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_694 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_210_1188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18164_ VGND VPWR _04077_ _03965_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15376_ VGND VPWR _00022_ _10837_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12588_ VPWR VGND VPWR VGND _08147_ keymem.key_mem\[6\]\[43\] _07739_ keymem.key_mem\[2\]\[43\]
+ _07698_ _08148_ sky130_fd_sc_hd__a221o_2
XFILLER_0_182_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_262_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14327_ VPWR VGND VGND VPWR _09053_ _09797_ _09056_ sky130_fd_sc_hd__nor2_2
X_17115_ VPWR VGND VGND VPWR _10732_ _03230_ key[69] sky130_fd_sc_hd__nor2_2
X_18095_ VPWR VGND VPWR VGND _04014_ _04010_ _04013_ sky130_fd_sc_hd__or2_2
XFILLER_0_20_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17046_ _02831_ _03168_ keymem.prev_key1_reg\[62\] _02832_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_14258_ VPWR VGND VPWR VGND _09728_ _09727_ sky130_fd_sc_hd__inv_2
XFILLER_0_257_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_223_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_382 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1276 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13209_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[104\] _07561_ keymem.key_mem\[1\]\[104\]
+ _07557_ _08708_ sky130_fd_sc_hd__a22o_2
X_14189_ VPWR VGND VPWR VGND _09656_ _09659_ _09657_ _09655_ _09660_ sky130_fd_sc_hd__or4_2
XFILLER_0_0_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_976 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18997_ VPWR VGND _04828_ _04827_ enc_block.round_key\[57\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_225_626 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17948_ VGND VPWR VPWR VGND _03896_ _03895_ keymem.prev_key0_reg\[106\] _03897_ sky130_fd_sc_hd__mux2_2
XFILLER_0_256_1358 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17879_ VGND VPWR _00225_ _03849_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_45_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_139_1178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19618_ VGND VPWR VPWR VGND _05205_ _05037_ keymem.key_mem\[12\]\[102\] _05212_ sky130_fd_sc_hd__mux2_2
XFILLER_0_215_1022 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_1128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20890_ VPWR VGND keymem.key_mem\[7\]\[56\] _05890_ _05886_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_75_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19549_ VPWR VGND keymem.key_mem\[12\]\[69\] _05176_ _05173_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_7_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22560_ VGND VPWR VPWR VGND _06750_ keymem.key_mem\[1\]\[83\] _03356_ _06765_ sky130_fd_sc_hd__mux2_2
XFILLER_0_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21511_ VGND VPWR _01488_ _06218_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_812 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22491_ VGND VPWR _06736_ _03859_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_228_1416 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24230_ VGND VPWR VPWR VGND clk _00723_ reset_n keymem.key_mem\[11\]\[95\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_145_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21442_ VGND VPWR _01455_ _06182_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_9_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_17_889 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_86_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24161_ VGND VPWR VPWR VGND clk _00654_ reset_n keymem.key_mem\[11\]\[26\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_44_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21373_ VGND VPWR _01422_ _06146_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_1246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23112_ VGND VPWR VPWR VGND _07032_ _07034_ keymem.prev_key1_reg\[96\] _07035_ sky130_fd_sc_hd__mux2_2
X_20324_ VGND VPWR VPWR VGND _05580_ _03035_ keymem.key_mem\[9\]\[48\] _05588_ sky130_fd_sc_hd__mux2_2
XFILLER_0_222_1004 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_128_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24092_ VGND VPWR VPWR VGND clk _00585_ reset_n keymem.key_mem\[12\]\[85\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_226_1184 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_12_550 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_141_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_84_2_Right_156 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23043_ VGND VPWR VPWR VGND _06992_ _03233_ keymem.prev_key1_reg\[69\] _06993_ sky130_fd_sc_hd__mux2_2
X_20255_ VGND VPWR VPWR VGND _05546_ _11149_ keymem.key_mem\[9\]\[15\] _05552_ sky130_fd_sc_hd__mux2_2
XFILLER_0_256_751 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20186_ VGND VPWR _00868_ _05513_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_122_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_486 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24994_ VGND VPWR VPWR VGND clk _01487_ reset_n keymem.key_mem\[5\]\[91\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_255_294 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_157_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1211 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_118_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23945_ VGND VPWR VPWR VGND clk _00438_ reset_n keymem.key_mem\[13\]\[66\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_1222 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_262_Right_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11890_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[16\] dec_new_block\[112\]
+ _07509_ sky130_fd_sc_hd__mux2_2
X_23876_ VGND VPWR VPWR VGND clk _00369_ reset_n enc_block.block_w2_reg\[29\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25615_ VGND VPWR VPWR VGND clk _02108_ reset_n keymem.key_mem\[0\]\[72\] sky130_fd_sc_hd__dfrtp_2
X_22827_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[126\] _06839_ _03864_ _05087_ _02162_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_6_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13560_ VGND VPWR VPWR VGND _09031_ _09017_ _09008_ _09032_ sky130_fd_sc_hd__or3_2
X_25546_ VGND VPWR VPWR VGND clk _02039_ reset_n keymem.key_mem\[0\]\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_109_302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22758_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[74\] _06837_ _06836_ _04989_ _02110_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_109_324 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12511_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[36\] _07759_ keymem.key_mem\[8\]\[36\]
+ _07540_ _08078_ sky130_fd_sc_hd__a22o_2
X_21709_ VGND VPWR VPWR VGND _06319_ _03118_ keymem.key_mem\[4\]\[57\] _06324_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_33_Left_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13491_ VGND VPWR VGND VPWR _08963_ _08962_ _08961_ keymem.prev_key1_reg\[3\] _08956_
+ _08943_ sky130_fd_sc_hd__a32o_2
X_25477_ VGND VPWR VPWR VGND clk _01970_ reset_n keymem.key_mem\[1\]\[62\] sky130_fd_sc_hd__dfrtp_2
X_22689_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[33\] _06790_ _06789_ _04922_ _02069_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_168_1330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15230_ VPWR VGND VGND VPWR _10535_ _10693_ _10498_ sky130_fd_sc_hd__nor2_2
XFILLER_0_129_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24428_ VGND VPWR VPWR VGND clk _00921_ reset_n keymem.key_mem\[9\]\[37\] sky130_fd_sc_hd__dfrtp_2
X_12442_ VGND VPWR enc_block.round_key\[29\] _08015_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_168_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_34_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_69_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_129_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15161_ VGND VPWR VGND VPWR _10618_ _10563_ _10584_ _10574_ _10625_ sky130_fd_sc_hd__a31o_2
XFILLER_0_50_612 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12373_ VGND VPWR enc_block.round_key\[23\] _07952_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24359_ VGND VPWR VPWR VGND clk _00852_ reset_n keymem.key_mem\[10\]\[96\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_65_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14112_ VPWR VGND VGND VPWR _09440_ _09583_ _09582_ sky130_fd_sc_hd__nor2_2
XFILLER_0_22_336 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15092_ VPWR VGND VPWR VGND _10447_ _10466_ _10403_ _10392_ _10556_ sky130_fd_sc_hd__or4_2
XFILLER_0_10_509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_678 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_729 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18920_ VPWR VGND VPWR VGND _04758_ block[49] _04744_ enc_block.block_w3_reg\[17\]
+ _04666_ _04759_ sky130_fd_sc_hd__a221o_2
X_14043_ VGND VPWR VGND VPWR _09515_ keymem.round_ctr_reg\[0\] _08933_ keymem.round_ctr_reg\[1\]
+ sky130_fd_sc_hd__and3b_2
XFILLER_0_30_391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18851_ VGND VPWR VGND VPWR _04697_ _03982_ _04696_ _04695_ sky130_fd_sc_hd__o21a_2
XPHY_EDGE_ROW_42_Left_310 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1087 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17802_ VPWR VGND VPWR VGND _03137_ _03797_ keymem.prev_key0_reg\[59\] _03788_ _00200_
+ sky130_fd_sc_hd__a22o_2
X_18782_ VPWR VGND VPWR VGND _04634_ _04550_ _04633_ enc_block.block_w2_reg\[3\] _04602_
+ _00343_ sky130_fd_sc_hd__a221o_2
XFILLER_0_101_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15994_ VPWR VGND VPWR VGND _11449_ keymem.prev_key1_reg\[81\] sky130_fd_sc_hd__inv_2
X_17733_ VGND VPWR _00174_ _03754_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_13_Right_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14945_ VGND VPWR _10409_ _10408_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_76_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_136_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17664_ VGND VPWR VPWR VGND _03703_ _03705_ keymem.prev_key0_reg\[13\] _03706_ sky130_fd_sc_hd__mux2_2
XFILLER_0_37_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14876_ VPWR VGND VGND VPWR _09040_ _10341_ _09051_ sky130_fd_sc_hd__nor2_2
XFILLER_0_230_640 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_72_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19403_ VGND VPWR VGND VPWR _05097_ keymem.key_mem_we _09725_ _05093_ _00501_ sky130_fd_sc_hd__a31o_2
X_16615_ VPWR VGND _02771_ _02770_ keymem.prev_key0_reg\[124\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_13827_ VGND VPWR _09299_ _09298_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17595_ VPWR VGND VPWR VGND _03653_ _03650_ _03649_ key[253] _08929_ _03654_ sky130_fd_sc_hd__a221o_2
XFILLER_0_106_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19334_ VPWR VGND keymem.key_mem_we _05050_ _03543_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_174_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13758_ VPWR VGND VGND VPWR _09065_ _09230_ _09041_ sky130_fd_sc_hd__nor2_2
X_16546_ VGND VPWR _02705_ _02702_ _02704_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_130_1_Right_731 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_174_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_112_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12709_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[54\] _08145_ _08257_ _08251_ _08258_
+ sky130_fd_sc_hd__o22a_2
X_19265_ VGND VPWR VGND VPWR _05005_ keymem.key_mem_we _03356_ _04999_ _00455_ sky130_fd_sc_hd__a31o_2
X_13689_ VGND VPWR VGND VPWR _09148_ _09160_ _09090_ _09069_ _09161_ sky130_fd_sc_hd__o22a_2
X_16477_ VGND VPWR VGND VPWR _02637_ _02612_ _02638_ _09240_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_127_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18216_ VGND VPWR VGND VPWR _04125_ _03972_ _11018_ _10993_ sky130_fd_sc_hd__o21a_2
XFILLER_0_112_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15428_ VGND VPWR VGND VPWR _10885_ _10590_ _10886_ _10887_ _10889_ _10888_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_13_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Right_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19196_ VGND VPWR _00427_ _04964_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_198_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18147_ VPWR VGND VGND VPWR _04062_ _04004_ _11104_ sky130_fd_sc_hd__nand2_2
X_15359_ _10818_ _10821_ _10817_ _10819_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_198_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_83_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1362 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_48_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18078_ VGND VPWR _03998_ enc_block.block_w0_reg\[26\] _03997_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_262_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_257_526 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_22_881 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_40_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17029_ VGND VPWR _03152_ _09543_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_81_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20040_ VGND VPWR _00798_ _05437_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_123_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_570 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_225_423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_197_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_193_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21991_ VPWR VGND keymem.key_mem\[3\]\[59\] _06476_ _06469_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_154_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_319 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23730_ keymem.prev_key0_reg\[86\] clk _00227_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_256_1199 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_94_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20942_ VPWR VGND keymem.key_mem\[7\]\[80\] _05918_ _05899_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_55_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_459 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_234_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23661_ keymem.prev_key0_reg\[17\] clk _00158_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20873_ VGND VPWR VPWR VGND _05880_ _04950_ keymem.key_mem\[7\]\[48\] _05881_ sky130_fd_sc_hd__mux2_2
XFILLER_0_221_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25400_ VGND VPWR VPWR VGND clk _01893_ reset_n keymem.key_mem\[2\]\[113\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_7_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22612_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[122\] _06756_ _03793_ _05079_ _02030_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_113_1148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23592_ VGND VPWR VPWR VGND clk _00093_ reset_n keymem.key_mem\[14\]\[81\] sky130_fd_sc_hd__dfrtp_2
X_25331_ VGND VPWR VPWR VGND clk _01824_ reset_n keymem.key_mem\[2\]\[44\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_130_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22543_ VGND VPWR _01979_ _06759_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_40_Right_40 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25262_ VGND VPWR VPWR VGND clk _01755_ reset_n keymem.key_mem\[3\]\[103\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_165_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_45_962 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22474_ VGND VPWR _01938_ _06731_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_664 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_118_187 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_267_1284 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_601 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_60_910 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24213_ VGND VPWR VPWR VGND clk _00706_ reset_n keymem.key_mem\[11\]\[78\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_133_146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21425_ VGND VPWR VPWR VGND _06173_ _03067_ keymem.key_mem\[5\]\[51\] _06174_ sky130_fd_sc_hd__mux2_2
XFILLER_0_165_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25193_ VGND VPWR VPWR VGND clk _01686_ reset_n keymem.key_mem\[3\]\[34\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_206_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24144_ VGND VPWR VPWR VGND clk _00637_ reset_n keymem.key_mem\[11\]\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_976 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21356_ VGND VPWR _01414_ _06137_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_114_382 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20307_ VGND VPWR VPWR VGND _05569_ _02955_ keymem.key_mem\[9\]\[40\] _05579_ sky130_fd_sc_hd__mux2_2
XFILLER_0_206_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_202_1408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24075_ VGND VPWR VPWR VGND clk _00568_ reset_n keymem.key_mem\[12\]\[68\] sky130_fd_sc_hd__dfrtp_2
X_21287_ VGND VPWR VPWR VGND _06098_ _03585_ keymem.key_mem\[6\]\[115\] _06100_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_85_2_Right_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_203_Left_470 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23026_ VGND VPWR VPWR VGND _02239_ _03167_ _03171_ _06925_ _06982_ sky130_fd_sc_hd__o31a_2
X_20238_ VGND VPWR VPWR VGND _05535_ _10369_ keymem.key_mem\[9\]\[7\] _05543_ sky130_fd_sc_hd__mux2_2
XFILLER_0_204_1290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_102_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_217_924 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_592 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_243_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20169_ VGND VPWR VPWR VGND _05504_ _03518_ keymem.key_mem\[10\]\[104\] _05505_ sky130_fd_sc_hd__mux2_2
XFILLER_0_102_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_243_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12991_ VGND VPWR VGND VPWR _08016_ keymem.key_mem\[7\]\[82\] _08507_ _08509_ _08512_
+ _08511_ sky130_fd_sc_hd__a2111o_2
X_24977_ VGND VPWR VPWR VGND clk _01470_ reset_n keymem.key_mem\[5\]\[74\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_172_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14730_ VPWR VGND VGND VPWR _09122_ _10196_ _09095_ sky130_fd_sc_hd__nor2_2
X_11942_ VGND VPWR _07545_ _07544_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23928_ VGND VPWR VPWR VGND clk _00421_ reset_n keymem.key_mem\[13\]\[49\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_252_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14661_ VGND VPWR VPWR VGND _09335_ _09247_ _09332_ _10128_ sky130_fd_sc_hd__or3_2
X_11873_ VGND VPWR result[103] _07500_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23859_ VGND VPWR VPWR VGND clk _00352_ reset_n enc_block.block_w2_reg\[12\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_15_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16400_ VGND VPWR VPWR VGND _02561_ _02562_ _02558_ _02557_ _11236_ _11379_ sky130_fd_sc_hd__o2111ai_2
X_13612_ VPWR VGND VGND VPWR _09067_ _09080_ _09084_ _09083_ _09082_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_197_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14592_ VPWR VGND VPWR VGND _10060_ _09765_ _10059_ sky130_fd_sc_hd__or2_2
X_17380_ VGND VPWR VPWR VGND _03467_ keymem.key_mem\[14\]\[96\] _03466_ _03468_ sky130_fd_sc_hd__mux2_2
XFILLER_0_200_857 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_156_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13543_ VGND VPWR _09015_ _08997_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16331_ VPWR VGND VGND VPWR _02494_ _02490_ _02493_ sky130_fd_sc_hd__nand2_2
X_25529_ VGND VPWR VPWR VGND clk _02022_ reset_n keymem.key_mem\[1\]\[114\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_55_759 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_54_236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_207_Right_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16262_ VGND VPWR VGND VPWR _11527_ _11386_ _11284_ _11377_ _11422_ _02426_ sky130_fd_sc_hd__o32a_2
X_19050_ VPWR VGND VGND VPWR _04600_ _04875_ _04301_ sky130_fd_sc_hd__nor2_2
X_13474_ VPWR VGND VGND VPWR enc_block.block_w1_reg\[2\] enc_block.sword_ctr_reg\[0\]
+ _08946_ sky130_fd_sc_hd__or2b_2
XFILLER_0_168_1171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15213_ VPWR VGND VPWR VGND _10675_ _10676_ _10673_ _10674_ sky130_fd_sc_hd__or3b_2
X_18001_ VGND VPWR VGND VPWR _03730_ keymem.prev_key0_reg\[123\] _03932_ _03638_ _00264_
+ sky130_fd_sc_hd__a2bb2o_2
X_12425_ VPWR VGND VPWR VGND _07999_ keymem.key_mem\[14\]\[28\] _07583_ keymem.key_mem\[10\]\[28\]
+ _07561_ _08000_ sky130_fd_sc_hd__a221o_2
X_16193_ VPWR VGND VPWR VGND _02357_ _02358_ _11231_ _11595_ sky130_fd_sc_hd__or3b_2
XFILLER_0_246_1368 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15144_ VGND VPWR _10608_ _10411_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12356_ VPWR VGND VPWR VGND _07936_ keymem.key_mem\[3\]\[22\] _07651_ keymem.key_mem\[14\]\[22\]
+ _07744_ _07937_ sky130_fd_sc_hd__a221o_2
XFILLER_0_129_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_105_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_244_1081 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_239_526 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_168_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15075_ VGND VPWR VPWR VGND _10463_ _10464_ _10473_ _10539_ sky130_fd_sc_hd__or3_2
XFILLER_0_26_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19952_ VGND VPWR VPWR VGND _05389_ _09725_ keymem.key_mem\[10\]\[1\] _05391_ sky130_fd_sc_hd__mux2_2
XFILLER_0_10_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12287_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[17\] _07659_ keymem.key_mem\[7\]\[17\]
+ _07872_ _07873_ sky130_fd_sc_hd__a22o_2
X_14026_ VPWR VGND VGND VPWR _09487_ _09498_ _09401_ sky130_fd_sc_hd__nor2_2
X_18903_ VPWR VGND VPWR VGND _04743_ _04664_ _04742_ enc_block.block_w2_reg\[15\]
+ _04709_ _00355_ sky130_fd_sc_hd__a221o_2
XFILLER_0_208_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19883_ VGND VPWR VPWR VGND _05350_ keymem.key_mem\[11\]\[98\] _03480_ _05353_ sky130_fd_sc_hd__mux2_2
XFILLER_0_235_721 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_216_Right_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18834_ VGND VPWR VPWR VGND _04600_ enc_block.block_w2_reg\[8\] _04074_ _04682_ sky130_fd_sc_hd__mux2_2
XFILLER_0_93_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_765 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_207_456 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18765_ VPWR VGND VGND VPWR _04619_ _04615_ _04617_ sky130_fd_sc_hd__nand2_2
X_15977_ VPWR VGND VGND VPWR _11433_ _11241_ _11380_ sky130_fd_sc_hd__nand2_2
XFILLER_0_253_1317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17716_ VPWR VGND VGND VPWR _03743_ _03744_ _03731_ sky130_fd_sc_hd__nor2_2
XFILLER_0_165_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14928_ VGND VPWR VGND VPWR _10392_ _10391_ _10390_ keymem.prev_key1_reg\[9\] _08955_
+ _08942_ sky130_fd_sc_hd__a32o_2
X_18696_ VPWR VGND VPWR VGND _04556_ block[91] _04487_ enc_block.block_w1_reg\[27\]
+ _04543_ _04557_ sky130_fd_sc_hd__a221o_2
XFILLER_0_76_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_651 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17647_ VGND VPWR VPWR VGND _03691_ key[136] keymem.prev_key1_reg\[8\] _03694_ sky130_fd_sc_hd__mux2_2
X_14859_ VGND VPWR VPWR VGND keylen _10324_ _10323_ _10319_ _10318_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_37_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17578_ VPWR VGND VPWR VGND _03637_ _10323_ _03639_ _03638_ keylen sky130_fd_sc_hd__a211oi_2
XFILLER_0_42_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19317_ VGND VPWR _00474_ _05038_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_225_Right_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16529_ VGND VPWR _02689_ _02688_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_131_1_Right_732 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19248_ VPWR VGND keymem.key_mem_we _04995_ _03306_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_45_269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_147_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_612 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_118_1_Left_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19179_ VGND VPWR VPWR VGND _04951_ _04953_ keymem.key_mem\[13\]\[49\] _04954_ sky130_fd_sc_hd__mux2_2
XFILLER_0_147_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21210_ VGND VPWR _01346_ _06059_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_108_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22190_ VGND VPWR VPWR VGND _06578_ _02688_ keymem.key_mem\[2\]\[24\] _06582_ sky130_fd_sc_hd__mux2_2
XFILLER_0_48_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21141_ VGND VPWR _01313_ _06023_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_13_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_857 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_572 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21072_ VGND VPWR _01280_ _05987_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_257_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_160_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20023_ VGND VPWR _00790_ _05428_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24900_ VGND VPWR VPWR VGND clk _01393_ reset_n keymem.key_mem\[6\]\[125\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_540 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_226_765 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24831_ VGND VPWR VPWR VGND clk _01324_ reset_n keymem.key_mem\[6\]\[56\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_158_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_50 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24762_ VGND VPWR VPWR VGND clk _01255_ reset_n keymem.key_mem\[7\]\[115\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_158_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21974_ VGND VPWR VGND VPWR _06466_ keymem.key_mem_we _03068_ _06446_ _01703_ sky130_fd_sc_hd__a31o_2
XFILLER_0_119_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23713_ keymem.prev_key0_reg\[69\] clk _00210_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_234_1250 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20925_ VGND VPWR _01212_ _05908_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24693_ VGND VPWR VPWR VGND clk _01186_ reset_n keymem.key_mem\[7\]\[46\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_7_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23644_ keymem.prev_key0_reg\[0\] clk _00141_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20856_ VGND VPWR VPWR VGND _05867_ _04935_ keymem.key_mem\[7\]\[40\] _05872_ sky130_fd_sc_hd__mux2_2
XFILLER_0_95_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23575_ VGND VPWR VPWR VGND clk _00076_ reset_n keymem.key_mem\[14\]\[64\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_748 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20787_ VGND VPWR VGND VPWR _05834_ keymem.key_mem_we _10662_ _05821_ _01148_ sky130_fd_sc_hd__a31o_2
XFILLER_0_64_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25314_ VGND VPWR VPWR VGND clk _01807_ reset_n keymem.key_mem\[2\]\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_106_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22526_ VGND VPWR VPWR VGND _06750_ keymem.key_mem\[1\]\[63\] _03184_ _06751_ sky130_fd_sc_hd__mux2_2
XFILLER_0_228_1010 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_973 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_472 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_91_386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25245_ VGND VPWR VPWR VGND clk _01738_ reset_n keymem.key_mem\[3\]\[86\] sky130_fd_sc_hd__dfrtp_2
X_22457_ VGND VPWR _01930_ _06722_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12210_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[11\] _07582_ keymem.key_mem\[6\]\[11\]
+ _07564_ _07802_ sky130_fd_sc_hd__a22o_2
X_21408_ VGND VPWR VPWR VGND _06162_ _02985_ keymem.key_mem\[5\]\[43\] _06165_ sky130_fd_sc_hd__mux2_2
XFILLER_0_66_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13190_ VPWR VGND VPWR VGND keymem.key_mem\[4\]\[102\] _07550_ keymem.key_mem\[1\]\[102\]
+ _07556_ _08691_ sky130_fd_sc_hd__a22o_2
X_25176_ VGND VPWR VPWR VGND clk _01669_ reset_n keymem.key_mem\[3\]\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_199_91 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22388_ VGND VPWR _01898_ _06685_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_248_312 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24127_ VGND VPWR VPWR VGND clk _00620_ reset_n keymem.key_mem\[12\]\[120\] sky130_fd_sc_hd__dfrtp_2
X_12141_ VGND VPWR _07737_ _07558_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21339_ VGND VPWR VPWR VGND _06128_ _10835_ keymem.key_mem\[5\]\[10\] _06129_ sky130_fd_sc_hd__mux2_2
XFILLER_0_27_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24058_ VGND VPWR VPWR VGND clk _00551_ reset_n keymem.key_mem\[12\]\[51\] sky130_fd_sc_hd__dfrtp_2
X_12072_ VGND VPWR _07672_ _07592_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_86_2_Right_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15900_ VPWR VGND VGND VPWR _11174_ _11356_ _11263_ sky130_fd_sc_hd__nor2_2
X_23009_ VGND VPWR VPWR VGND _06960_ _06972_ keymem.prev_key1_reg\[55\] _06973_ sky130_fd_sc_hd__mux2_2
XFILLER_0_263_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_1084 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_8_Left_276 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16880_ VPWR VGND VPWR VGND _03017_ keymem.prev_key1_reg\[47\] sky130_fd_sc_hd__inv_2
XFILLER_0_21_1057 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15831_ VPWR VGND VGND VPWR _11287_ _11286_ _11221_ sky130_fd_sc_hd__nand2_2
XFILLER_0_176_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18550_ VPWR VGND _04426_ _04354_ enc_block.block_w0_reg\[4\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15762_ VGND VPWR _11218_ _11217_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12974_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[81\] _07779_ keymem.key_mem\[6\]\[81\]
+ _07657_ _08496_ sky130_fd_sc_hd__a22o_2
XFILLER_0_235_1047 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_73_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17501_ VGND VPWR VGND VPWR _03571_ _09637_ _03570_ _03569_ _03572_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_137_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14713_ VPWR VGND VGND VPWR _09114_ _10180_ _09658_ sky130_fd_sc_hd__nor2_2
X_18481_ VPWR VGND _04364_ enc_block.block_w1_reg\[29\] enc_block.block_w1_reg\[28\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_217_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11925_ VGND VPWR VPWR VGND encdec enc_block.round\[3\] dec_round_nr\[3\] _07528_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_86_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_234_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15693_ VGND VPWR VPWR VGND _11041_ keymem.key_mem\[14\]\[15\] _11149_ _11150_ sky130_fd_sc_hd__mux2_2
XFILLER_0_34_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1394 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17432_ VGND VPWR _00115_ _03512_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_213_1345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14644_ VGND VPWR VGND VPWR _09400_ _09418_ _09354_ _09452_ _10111_ sky130_fd_sc_hd__o22a_2
X_11856_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[31\] dec_new_block\[95\]
+ _07492_ sky130_fd_sc_hd__mux2_2
X_14575_ VGND VPWR _10042_ _09302_ _10043_ _09350_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_17363_ VGND VPWR VPWR VGND _03384_ keymem.key_mem\[14\]\[94\] _03452_ _03453_ sky130_fd_sc_hd__mux2_2
XFILLER_0_27_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11787_ VGND VPWR result[60] _07457_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_248_1419 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_250_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19102_ VPWR VGND keymem.key_mem\[13\]\[20\] _04906_ _04903_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16314_ VPWR VGND VPWR VGND _02475_ _02469_ _02478_ _02477_ keylen sky130_fd_sc_hd__a211oi_2
X_13526_ VPWR VGND VPWR VGND _08982_ _08997_ _08991_ _08977_ _08998_ sky130_fd_sc_hd__or4_2
X_17294_ VGND VPWR VPWR VGND _03389_ _02947_ _03391_ _09514_ _03390_ sky130_fd_sc_hd__o211a_2
XFILLER_0_250_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_148_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19033_ VGND VPWR VGND VPWR _04859_ _04266_ _04600_ _04860_ enc_block.block_w2_reg\[29\]
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_152_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13457_ VGND VPWR _08929_ _08928_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16245_ VGND VPWR _02410_ _02409_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_42_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_148_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12408_ VGND VPWR _07984_ _07583_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_2_325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_976 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_258_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_152_285 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_84_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13388_ VPWR VGND VPWR VGND _08868_ keymem.key_mem\[14\]\[122\] _08032_ keymem.key_mem\[6\]\[122\]
+ _07771_ _08869_ sky130_fd_sc_hd__a221o_2
X_16176_ VGND VPWR _00030_ _02341_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_45_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15127_ _10590_ _10591_ _10463_ _10487_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_12339_ VGND VPWR VGND VPWR _07922_ _07648_ keymem.key_mem\[2\]\[20\] _07917_ _07921_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_10_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_224_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15058_ VGND VPWR _10522_ _10521_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_266_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19935_ VGND VPWR VPWR VGND _05372_ keymem.key_mem\[11\]\[123\] _03640_ _05380_ sky130_fd_sc_hd__mux2_2
XFILLER_0_254_304 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_195_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_259_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14009_ VPWR VGND VGND VPWR _09437_ _09323_ _09481_ _09479_ _09480_ _09478_ sky130_fd_sc_hd__o32ai_2
XFILLER_0_248_890 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_103_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19866_ VGND VPWR VPWR VGND _05339_ keymem.key_mem\[11\]\[90\] _03418_ _05344_ sky130_fd_sc_hd__mux2_2
X_18817_ VGND VPWR _04666_ _03977_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19797_ VGND VPWR VPWR VGND _05303_ keymem.key_mem\[11\]\[57\] _03119_ _05308_ sky130_fd_sc_hd__mux2_2
XFILLER_0_155_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18748_ VGND VPWR _04603_ enc_block.block_w1_reg\[0\] enc_block.block_w1_reg\[7\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_231_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18679_ VPWR VGND VGND VPWR _04512_ _04542_ _04248_ sky130_fd_sc_hd__nor2_2
XFILLER_0_235_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_144_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_203_481 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_77_147 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20710_ VGND VPWR VPWR VGND _05783_ _03511_ keymem.key_mem\[8\]\[103\] _05791_ sky130_fd_sc_hd__mux2_2
XFILLER_0_77_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21690_ VGND VPWR VPWR VGND _06308_ _03035_ keymem.key_mem\[4\]\[48\] _06314_ sky130_fd_sc_hd__mux2_2
XFILLER_0_8_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20641_ VGND VPWR VPWR VGND _05747_ _03245_ keymem.key_mem\[8\]\[70\] _05755_ sky130_fd_sc_hd__mux2_2
XFILLER_0_50_1242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23360_ VPWR VGND VPWR VGND _07235_ block[15] _04837_ enc_block.block_w1_reg\[15\]
+ _04504_ _07236_ sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_132_1_Right_733 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20572_ VGND VPWR VPWR VGND _05714_ _02923_ keymem.key_mem\[8\]\[37\] _05719_ sky130_fd_sc_hd__mux2_2
XFILLER_0_50_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22311_ VGND VPWR VPWR VGND _06634_ _03346_ keymem.key_mem\[2\]\[82\] _06645_ sky130_fd_sc_hd__mux2_2
XFILLER_0_15_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23291_ VGND VPWR VPWR VGND _07093_ enc_block.block_w3_reg\[8\] _04074_ _07174_ sky130_fd_sc_hd__mux2_2
XFILLER_0_6_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25030_ VGND VPWR VPWR VGND clk _01523_ reset_n keymem.key_mem\[5\]\[127\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_143_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22242_ VGND VPWR VPWR VGND _06600_ _03046_ keymem.key_mem\[2\]\[49\] _06609_ sky130_fd_sc_hd__mux2_2
XFILLER_0_44_1002 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22173_ VGND VPWR VPWR VGND _06565_ _11446_ keymem.key_mem\[2\]\[16\] _06573_ sky130_fd_sc_hd__mux2_2
XFILLER_0_203_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21124_ VGND VPWR _01305_ _06014_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_160_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_258_1014 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_61_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21055_ VGND VPWR VPWR VGND _05972_ _10193_ keymem.key_mem\[6\]\[5\] _05978_ sky130_fd_sc_hd__mux2_2
XFILLER_0_219_1009 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20006_ VGND VPWR _00782_ _05419_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_198_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24814_ VGND VPWR VPWR VGND clk _01307_ reset_n keymem.key_mem\[6\]\[39\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_214_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_234 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25794_ keymem.prev_key1_reg\[110\] clk _02287_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_24745_ VGND VPWR VPWR VGND clk _01238_ reset_n keymem.key_mem\[7\]\[98\] sky130_fd_sc_hd__dfrtp_2
X_21957_ VGND VPWR _01695_ _06457_ VPWR VGND sky130_fd_sc_hd__buf_1
X_11710_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[22\] dec_new_block\[22\]
+ _07419_ sky130_fd_sc_hd__mux2_2
X_20908_ VPWR VGND keymem.key_mem\[7\]\[64\] _05900_ _05899_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_178_171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_56_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12690_ VPWR VGND VPWR VGND keymem.key_mem\[8\]\[53\] _07958_ keymem.key_mem\[1\]\[53\]
+ _07901_ _08240_ sky130_fd_sc_hd__a22o_2
X_24676_ VGND VPWR VPWR VGND clk _01169_ reset_n keymem.key_mem\[7\]\[29\] sky130_fd_sc_hd__dfrtp_2
X_21888_ VGND VPWR _06420_ _06403_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_166_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23627_ VGND VPWR VPWR VGND clk _00128_ reset_n keymem.key_mem\[14\]\[116\] sky130_fd_sc_hd__dfrtp_2
X_11641_ VGND VPWR VPWR VGND enc_block.round\[1\] enc_block.round\[2\] _07380_ enc_block.round\[3\]
+ _07379_ sky130_fd_sc_hd__o211a_2
X_20839_ VGND VPWR _01172_ _05862_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_210_996 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_132_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_193_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14360_ VGND VPWR VGND VPWR _09148_ _09083_ _09036_ _09203_ _09830_ sky130_fd_sc_hd__o22a_2
XFILLER_0_64_342 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23558_ VGND VPWR VPWR VGND clk _00059_ reset_n keymem.key_mem\[14\]\[47\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_25_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13311_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[114\] _08391_ keymem.key_mem\[6\]\[114\]
+ _07656_ _08800_ sky130_fd_sc_hd__a22o_2
X_22509_ VGND VPWR _01962_ _06742_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14291_ VPWR VGND VGND VPWR _09343_ _09366_ _09761_ _09450_ _09495_ sky130_fd_sc_hd__o22ai_2
X_23489_ VGND VPWR _07350_ enc_block.block_w0_reg\[21\] enc_block.block_w0_reg\[22\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_16030_ VPWR VGND VPWR VGND _11485_ _11483_ _11484_ sky130_fd_sc_hd__or2_2
X_13242_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[107\] _07725_ keymem.key_mem\[14\]\[107\]
+ _07666_ _08738_ sky130_fd_sc_hd__a22o_2
XFILLER_0_243_1338 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25228_ VGND VPWR VPWR VGND clk _01721_ reset_n keymem.key_mem\[3\]\[69\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_773 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_27_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13173_ VGND VPWR VGND VPWR _07542_ keymem.key_mem\[8\]\[100\] _08672_ _08673_ _08676_
+ _08675_ sky130_fd_sc_hd__a2111o_2
X_25159_ VGND VPWR VPWR VGND clk _01652_ reset_n keymem.key_mem\[3\]\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_676 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12124_ VGND VPWR _07721_ _07706_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17981_ VGND VPWR VPWR VGND _03281_ key[245] keymem.prev_key1_reg\[117\] _03919_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_102_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19720_ VGND VPWR _00648_ _05267_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16932_ VGND VPWR VPWR VGND _03065_ _02403_ _09866_ _03064_ _09533_ sky130_fd_sc_hd__o31ai_2
X_12055_ VGND VPWR _07655_ _07654_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_87_2_Right_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_263_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19651_ VGND VPWR _00617_ _05229_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16863_ VPWR VGND VPWR VGND _03002_ keymem.prev_key1_reg\[45\] sky130_fd_sc_hd__inv_2
XFILLER_0_245_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_254_1412 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18602_ VGND VPWR VGND VPWR _04472_ _04470_ _04473_ _03965_ sky130_fd_sc_hd__a21oi_2
X_15814_ VGND VPWR _11270_ _11269_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19582_ VGND VPWR _00584_ _05193_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_204_234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_232_554 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16794_ VGND VPWR VPWR VGND _02936_ _10329_ _02939_ _02938_ _02937_ sky130_fd_sc_hd__o211a_2
XFILLER_0_172_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18533_ VGND VPWR _04411_ _04409_ _04410_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_245_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15745_ VPWR VGND VPWR VGND _11201_ enc_block.block_w0_reg\[21\] _08995_ sky130_fd_sc_hd__or2_2
X_12957_ VGND VPWR VGND VPWR _07780_ keymem.key_mem\[5\]\[79\] _08477_ _08479_ _08481_
+ _08480_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_38_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11908_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[25\] dec_new_block\[121\]
+ _07518_ sky130_fd_sc_hd__mux2_2
X_18464_ VGND VPWR _04349_ enc_block.round_key\[67\] _04348_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_213_1142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15676_ VGND VPWR VGND VPWR _10516_ _10682_ _10639_ _11133_ sky130_fd_sc_hd__a21o_2
XFILLER_0_59_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12888_ VPWR VGND VPWR VGND _08418_ keymem.key_mem\[5\]\[72\] _07597_ keymem.key_mem\[4\]\[72\]
+ _07552_ _08419_ sky130_fd_sc_hd__a221o_2
XFILLER_0_150_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_157_344 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17415_ VPWR VGND VGND VPWR _03498_ _09534_ _03497_ sky130_fd_sc_hd__nand2_2
XFILLER_0_261_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_184_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14627_ VGND VPWR _10094_ _10092_ _10095_ _10089_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_11839_ VGND VPWR result[86] _07483_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18395_ VPWR VGND VGND VPWR _04287_ _04044_ _04285_ sky130_fd_sc_hd__nand2_2
XFILLER_0_172_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_150_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_128_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17346_ VGND VPWR VGND VPWR _02804_ _02803_ _02708_ _03437_ sky130_fd_sc_hd__a21o_2
X_14558_ VPWR VGND VPWR VGND _09828_ _10025_ _10024_ _10023_ _10026_ sky130_fd_sc_hd__or4_2
XFILLER_0_28_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_537 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13509_ VPWR VGND VPWR VGND _08981_ enc_block.block_w0_reg\[6\] _08952_ sky130_fd_sc_hd__or2_2
X_17277_ VGND VPWR _00097_ _03375_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14489_ VPWR VGND VGND VPWR _09089_ _08972_ _09958_ _09140_ _09124_ sky130_fd_sc_hd__o22ai_2
X_19016_ VPWR VGND VGND VPWR _04778_ _04845_ _04258_ sky130_fd_sc_hd__nor2_2
XFILLER_0_109_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16228_ VGND VPWR VGND VPWR _02377_ _02392_ _02393_ _02373_ _02382_ sky130_fd_sc_hd__nor4_2
XFILLER_0_130_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_261_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_23_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_109_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16159_ VPWR VGND VGND VPWR _11210_ _11313_ _11613_ _11218_ _11344_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_51_592 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_456 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_255_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_267_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_228_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_259_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19918_ VGND VPWR VPWR VGND _05361_ keymem.key_mem\[11\]\[115\] _03585_ _05371_ sky130_fd_sc_hd__mux2_2
XFILLER_0_255_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19849_ VGND VPWR VPWR VGND _05328_ keymem.key_mem\[11\]\[82\] _03347_ _05335_ sky130_fd_sc_hd__mux2_2
XFILLER_0_190_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22860_ VGND VPWR VPWR VGND _06878_ _09535_ keymem.prev_key1_reg\[0\] _06879_ sky130_fd_sc_hd__mux2_2
XFILLER_0_218_1064 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21811_ VGND VPWR _06377_ _06258_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22791_ VGND VPWR VPWR VGND _06784_ keymem.key_mem\[0\]\[95\] _03460_ _06856_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1278 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24530_ VGND VPWR VPWR VGND clk _01023_ reset_n keymem.key_mem\[8\]\[11\] sky130_fd_sc_hd__dfrtp_2
X_21742_ VGND VPWR VPWR VGND _06330_ _03267_ keymem.key_mem\[4\]\[73\] _06341_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24461_ VGND VPWR VPWR VGND clk _00954_ reset_n keymem.key_mem\[9\]\[70\] sky130_fd_sc_hd__dfrtp_2
X_21673_ VGND VPWR VPWR VGND _06297_ _02955_ keymem.key_mem\[4\]\[40\] _06305_ sky130_fd_sc_hd__mux2_2
XFILLER_0_11_1001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23412_ VPWR VGND VPWR VGND _07282_ _03950_ _07281_ enc_block.block_w3_reg\[20\]
+ _07126_ _02325_ sky130_fd_sc_hd__a221o_2
X_20624_ VGND VPWR VPWR VGND _05736_ _03172_ keymem.key_mem\[8\]\[62\] _05746_ sky130_fd_sc_hd__mux2_2
X_24392_ VGND VPWR VPWR VGND clk _00885_ reset_n keymem.key_mem\[9\]\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_11_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23343_ VGND VPWR VPWR VGND _07093_ enc_block.block_w3_reg\[13\] _07220_ _07221_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_62_846 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_133_1_Right_734 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20555_ VGND VPWR VPWR VGND _05703_ _02811_ keymem.key_mem\[8\]\[29\] _05710_ sky130_fd_sc_hd__mux2_2
XFILLER_0_149_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23274_ VPWR VGND _07158_ enc_block.block_w1_reg\[15\] enc_block.block_w2_reg\[6\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_61_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20486_ VGND VPWR _01009_ _05672_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25013_ VGND VPWR VPWR VGND clk _01506_ reset_n keymem.key_mem\[5\]\[110\] sky130_fd_sc_hd__dfrtp_2
X_22225_ VGND VPWR _06600_ _06553_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_225_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_827 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22156_ VGND VPWR _01788_ _06563_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_98_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21107_ VGND VPWR _01297_ _06005_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_22_1141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22087_ VGND VPWR VPWR VGND _06516_ _05043_ keymem.key_mem\[3\]\[105\] _06526_ sky130_fd_sc_hd__mux2_2
XFILLER_0_238_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21038_ VGND VPWR _01266_ _05967_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_22_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13860_ VGND VPWR VPWR VGND _09331_ _09315_ _09303_ _09332_ sky130_fd_sc_hd__or3_2
XFILLER_0_138_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12811_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[64\] _07536_ _08349_ _08345_ enc_block.round_key\[64\]
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_35_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13791_ enc_block.sword_ctr_reg\[1\] _09263_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[25\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_22989_ VGND VPWR _02223_ _06961_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25777_ keymem.prev_key1_reg\[93\] clk _02270_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_9_1057 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15530_ VPWR VGND VGND VPWR _10593_ _10989_ _10485_ sky130_fd_sc_hd__nor2_2
XFILLER_0_139_311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24728_ VGND VPWR VPWR VGND clk _01221_ reset_n keymem.key_mem\[7\]\[81\] sky130_fd_sc_hd__dfrtp_2
X_12742_ VGND VPWR enc_block.round_key\[57\] _08287_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_56_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15461_ VPWR VGND VGND VPWR _10644_ _10921_ _10667_ sky130_fd_sc_hd__nor2_2
X_12673_ VGND VPWR VGND VPWR _07808_ keymem.key_mem\[12\]\[51\] _08222_ _08224_ _08225_
+ _08069_ sky130_fd_sc_hd__a2111o_2
X_24659_ VGND VPWR VPWR VGND clk _01152_ reset_n keymem.key_mem\[7\]\[12\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_249_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17200_ VGND VPWR VPWR VGND _03296_ keymem.key_mem\[14\]\[77\] _03306_ _03307_ sky130_fd_sc_hd__mux2_2
XFILLER_0_139_388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14412_ VPWR VGND VPWR VGND _09880_ _09573_ _09879_ _09463_ _09496_ _09881_ sky130_fd_sc_hd__a221o_2
XFILLER_0_132_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_325 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18180_ VPWR VGND VGND VPWR _04091_ _04092_ _04077_ sky130_fd_sc_hd__nor2_2
X_15392_ VGND VPWR VGND VPWR _10496_ _10518_ _10411_ _10618_ _10853_ sky130_fd_sc_hd__o22a_2
XFILLER_0_71_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_249_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17131_ VPWR VGND VPWR VGND _03244_ _03242_ _03241_ key[198] _03027_ _03245_ sky130_fd_sc_hd__a221o_2
X_14343_ VPWR VGND VGND VPWR _09134_ _09813_ _09157_ sky130_fd_sc_hd__nor2_2
XFILLER_0_181_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14274_ VGND VPWR VGND VPWR _09380_ _09403_ _09426_ _09743_ _09744_ sky130_fd_sc_hd__o22a_2
X_17062_ VGND VPWR VGND VPWR _03183_ _03152_ key[191] _03177_ _03182_ sky130_fd_sc_hd__a211o_2
XFILLER_0_107_296 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_184_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_69_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16013_ VGND VPWR VGND VPWR _11467_ _11263_ _11377_ _11417_ _11468_ sky130_fd_sc_hd__a31o_2
XFILLER_0_61_890 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13225_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[105\] _08714_ _08722_ _08718_ _08723_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_122_266 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_58 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13156_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[99\] _07834_ keymem.key_mem\[8\]\[99\]
+ _08211_ _08660_ sky130_fd_sc_hd__a22o_2
XFILLER_0_209_315 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1291 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12107_ VGND VPWR _07705_ _07612_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_236_123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17964_ VGND VPWR _00252_ _03907_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13087_ VPWR VGND VPWR VGND _08597_ keymem.key_mem\[12\]\[92\] _07807_ keymem.key_mem\[8\]\[92\]
+ _07929_ _08598_ sky130_fd_sc_hd__a221o_2
XFILLER_0_236_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_104_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_264_465 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19703_ VGND VPWR _00640_ _05258_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16915_ VGND VPWR _02866_ key[50] _03049_ _10189_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_12038_ VGND VPWR _07639_ _07563_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_40_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_498 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17895_ VGND VPWR VGND VPWR _03792_ _02711_ _03727_ _03859_ _03861_ _03860_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_18_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_532 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19634_ VGND VPWR _00609_ _05220_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16846_ VGND VPWR VPWR VGND _02986_ keymem.key_mem\[14\]\[43\] _02985_ _02987_ sky130_fd_sc_hd__mux2_2
XFILLER_0_75_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_127_1_Left_394 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19565_ VGND VPWR _00576_ _05184_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_219_1395 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16777_ VGND VPWR _02924_ _02923_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_149_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13989_ VGND VPWR VGND VPWR _09423_ _09399_ _09461_ _09294_ sky130_fd_sc_hd__a21oi_2
X_18516_ _04394_ _04396_ _04065_ _04395_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_245_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15728_ VGND VPWR VGND VPWR _11184_ enc_block.sword_ctr_reg\[0\] enc_block.block_w1_reg\[23\]
+ enc_block.sword_ctr_reg\[1\] sky130_fd_sc_hd__and3b_2
X_19496_ VGND VPWR _00544_ _05147_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_34_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18447_ VGND VPWR _04333_ enc_block.block_w1_reg\[25\] _04332_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_157_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_150_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15659_ VPWR VGND VPWR VGND _10802_ _10863_ _10804_ _10781_ _11116_ sky130_fd_sc_hd__or4_2
XFILLER_0_111_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1002 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_51_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18378_ VPWR VGND VPWR VGND _04271_ block[124] _04213_ enc_block.block_w0_reg\[28\]
+ _04171_ _04272_ sky130_fd_sc_hd__a221o_2
XFILLER_0_50_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_846 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17329_ VGND VPWR VGND VPWR key[91] _09930_ _03421_ _03420_ _03422_ sky130_fd_sc_hd__o22a_2
XFILLER_0_50_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_70_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20340_ VGND VPWR _00939_ _05596_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_82_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_86_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_976 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_12_721 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_226_1366 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1257 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_45_1130 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20271_ VGND VPWR _00906_ _05560_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22010_ VPWR VGND VGND VPWR _06486_ keymem.key_mem\[3\]\[68\] _06406_ sky130_fd_sc_hd__nand2_2
XFILLER_0_122_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_243_Right_112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_255_443 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_122_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23961_ VGND VPWR VPWR VGND clk _00454_ reset_n keymem.key_mem\[13\]\[82\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_227_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25700_ keymem.prev_key1_reg\[16\] clk _02193_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_93_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22912_ VGND VPWR VGND VPWR _02195_ _06912_ _06882_ keymem.prev_key1_reg\[18\] sky130_fd_sc_hd__o21a_2
X_23892_ VGND VPWR VPWR VGND clk _00385_ reset_n keymem.key_mem\[13\]\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25631_ VGND VPWR VPWR VGND clk _02124_ reset_n keymem.key_mem\[0\]\[88\] sky130_fd_sc_hd__dfrtp_2
X_22843_ VGND VPWR VGND VPWR _02168_ _06870_ _06869_ keymem.rcon_logic.tmp_rcon\[5\]
+ _06867_ _06864_ sky130_fd_sc_hd__a32o_2
XFILLER_0_78_231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_195_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22774_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[85\] _06837_ _06836_ _05008_ _02121_
+ sky130_fd_sc_hd__a22o_2
X_25562_ VGND VPWR VPWR VGND clk _02055_ reset_n keymem.key_mem\[0\]\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21725_ VGND VPWR _01588_ _06332_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24513_ VGND VPWR VPWR VGND clk _01006_ reset_n keymem.key_mem\[9\]\[122\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_148_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_133_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25493_ VGND VPWR VPWR VGND clk _01986_ reset_n keymem.key_mem\[1\]\[78\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_136_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_802 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24444_ VGND VPWR VPWR VGND clk _00937_ reset_n keymem.key_mem\[9\]\[53\] sky130_fd_sc_hd__dfrtp_2
X_21656_ VGND VPWR VPWR VGND _06286_ _02873_ keymem.key_mem\[4\]\[32\] _06296_ sky130_fd_sc_hd__mux2_2
XFILLER_0_163_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_47_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_34_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_89_2_Left_560 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20607_ VGND VPWR _01065_ _05737_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24375_ VGND VPWR VPWR VGND clk _00868_ reset_n keymem.key_mem\[10\]\[112\] sky130_fd_sc_hd__dfrtp_2
X_21587_ VGND VPWR _06259_ _06258_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_34_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23326_ VGND VPWR _07205_ _07131_ _07204_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_144_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_827 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_134_1_Right_735 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_201_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20538_ VGND VPWR VPWR VGND _05692_ _02549_ keymem.key_mem\[8\]\[21\] _05701_ sky130_fd_sc_hd__mux2_2
XFILLER_0_104_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23257_ VGND VPWR _07143_ _07140_ _07142_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_244_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20469_ VGND VPWR VPWR VGND _05660_ _03600_ keymem.key_mem\[9\]\[117\] _05664_ sky130_fd_sc_hd__mux2_2
X_13010_ VPWR VGND VPWR VGND _08528_ keymem.key_mem\[13\]\[84\] _07730_ keymem.key_mem\[10\]\[84\]
+ _07743_ _08529_ sky130_fd_sc_hd__a221o_2
XFILLER_0_259_771 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22208_ VGND VPWR _01812_ _06591_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23188_ VGND VPWR _02302_ _07081_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_140_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22139_ VGND VPWR VPWR VGND _06554_ _09536_ keymem.key_mem\[2\]\[0\] _06555_ sky130_fd_sc_hd__mux2_2
XFILLER_0_101_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_219_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_140_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_192_1_Left_459 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_262_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_206_318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14961_ enc_block.sword_ctr_reg\[1\] _10425_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[14\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_101_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_262_969 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16700_ VGND VPWR VGND VPWR _02844_ keymem.prev_key1_reg\[127\] _02853_ _02843_ sky130_fd_sc_hd__nand3_2
X_13912_ VGND VPWR VGND VPWR _09378_ _09381_ _09294_ _09383_ _09384_ sky130_fd_sc_hd__o22a_2
X_17680_ VGND VPWR _00159_ _03716_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14892_ VPWR VGND VPWR VGND _10353_ _10356_ _10357_ _09642_ _10352_ sky130_fd_sc_hd__or4b_2
X_16631_ VGND VPWR _02787_ _02786_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13843_ VGND VPWR _09315_ _09314_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25829_ VGND VPWR VPWR VGND clk _02322_ reset_n enc_block.block_w3_reg\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_18_1029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_1078 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_251_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_916 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19350_ VGND VPWR VPWR VGND _05046_ _05060_ keymem.key_mem\[13\]\[113\] _05061_ sky130_fd_sc_hd__mux2_2
X_16562_ VGND VPWR _02721_ _02720_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13774_ VGND VPWR _09246_ _09245_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18301_ VPWR VGND VPWR VGND _04202_ _04189_ _04200_ enc_block.block_w0_reg\[20\]
+ _04097_ _00294_ sky130_fd_sc_hd__a221o_2
XFILLER_0_214_1270 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15513_ VGND VPWR _10972_ _10967_ _10973_ _10969_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_19281_ VGND VPWR VPWR VGND _04993_ _05015_ keymem.key_mem\[13\]\[89\] _05016_ sky130_fd_sc_hd__mux2_2
X_12725_ VPWR VGND VPWR VGND _08271_ keymem.key_mem\[4\]\[56\] _07914_ keymem.key_mem\[2\]\[56\]
+ _07698_ _08272_ sky130_fd_sc_hd__a221o_2
XFILLER_0_151_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16493_ VGND VPWR VGND VPWR _02652_ _02651_ _02654_ _02653_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_242_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18232_ VGND VPWR _04139_ _03957_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_112_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15444_ VPWR VGND VPWR VGND _10905_ keymem.prev_key1_reg\[75\] sky130_fd_sc_hd__inv_2
XFILLER_0_26_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12656_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[49\] _08145_ _08209_ _08205_ _08210_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_26_846 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18163_ VGND VPWR _04076_ _03979_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_5_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12587_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[43\] _07806_ keymem.key_mem\[4\]\[43\]
+ _07913_ _08147_ sky130_fd_sc_hd__a22o_2
X_15375_ VGND VPWR VPWR VGND _09864_ keymem.key_mem\[14\]\[10\] _10836_ _10837_ sky130_fd_sc_hd__mux2_2
XFILLER_0_0_1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_154_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17114_ VGND VPWR VPWR VGND _09717_ _10187_ keymem.prev_key0_reg\[69\] _03229_ sky130_fd_sc_hd__or3_2
X_14326_ VGND VPWR _09796_ _09795_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_40_304 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18094_ VGND VPWR _04013_ _04011_ _04012_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_262_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_52_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17045_ VGND VPWR VPWR VGND _09796_ key[62] _03167_ _03166_ _09931_ sky130_fd_sc_hd__o211a_2
XFILLER_0_64_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14257_ VPWR VGND _09727_ keymem.prev_key1_reg\[34\] keymem.prev_key1_reg\[2\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_262_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13208_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[104\] _07760_ keymem.key_mem\[4\]\[104\]
+ _07552_ _08707_ sky130_fd_sc_hd__a22o_2
XFILLER_0_150_394 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_110_236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14188_ VGND VPWR VGND VPWR _09159_ _09658_ _09659_ _09082_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_443 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13139_ VGND VPWR VGND VPWR _07842_ keymem.key_mem\[9\]\[97\] _08642_ _08644_ _08645_
+ _08599_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_195_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18996_ VPWR VGND VPWR VGND _04826_ block[57] _04744_ enc_block.block_w2_reg\[25\]
+ _04798_ _04827_ sky130_fd_sc_hd__a221o_2
X_17947_ VGND VPWR _03896_ _03673_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_40_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_249_Left_516 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_252_457 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17878_ VGND VPWR VPWR VGND _03836_ _03848_ keymem.prev_key0_reg\[84\] _03849_ sky130_fd_sc_hd__mux2_2
XFILLER_0_75_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19617_ VGND VPWR _00601_ _05211_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16829_ VGND VPWR VGND VPWR keylen _02971_ _02970_ _10323_ _10828_ _02968_ sky130_fd_sc_hd__a311oi_2
XFILLER_0_215_1034 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_18_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19548_ VGND VPWR VPWR VGND _00568_ _05095_ _03226_ _08922_ _05175_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_215_1078 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19479_ VGND VPWR VPWR VGND _05138_ _04927_ keymem.key_mem\[12\]\[36\] _05139_ sky130_fd_sc_hd__mux2_2
XFILLER_0_61_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21510_ VGND VPWR VPWR VGND _06209_ _03434_ keymem.key_mem\[5\]\[92\] _06218_ sky130_fd_sc_hd__mux2_2
XFILLER_0_8_545 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22490_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[42\] _06707_ _06706_ _04939_ _01950_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_56_470 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_835 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21441_ VGND VPWR VPWR VGND _06173_ _03139_ keymem.key_mem\[5\]\[59\] _06182_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_258_Left_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24160_ VGND VPWR VPWR VGND clk _00653_ reset_n keymem.key_mem\[11\]\[25\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_86_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21372_ VGND VPWR VPWR VGND _06140_ _02742_ keymem.key_mem\[5\]\[26\] _06146_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23111_ VGND VPWR VGND VPWR _03462_ _06928_ _03465_ _07034_ sky130_fd_sc_hd__a21o_2
X_20323_ VGND VPWR _00931_ _05587_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_1258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24091_ VGND VPWR VPWR VGND clk _00584_ reset_n keymem.key_mem\[12\]\[84\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_101_203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_90 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_101_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23042_ VGND VPWR _06992_ _06880_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_12_562 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_922 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20254_ VGND VPWR _00898_ _05551_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_101_258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_177_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_229_966 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_200_1325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20185_ VGND VPWR VPWR VGND _05504_ _03567_ keymem.key_mem\[10\]\[112\] _05513_ sky130_fd_sc_hd__mux2_2
XFILLER_0_86_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_239_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_267_Left_534 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_215_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24993_ VGND VPWR VPWR VGND clk _01486_ reset_n keymem.key_mem\[5\]\[90\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_157_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23944_ VGND VPWR VPWR VGND clk _00437_ reset_n keymem.key_mem\[13\]\[65\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_118_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_1234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_212_822 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_98_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1218 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23875_ VGND VPWR VPWR VGND clk _00368_ reset_n enc_block.block_w2_reg\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25614_ VGND VPWR VPWR VGND clk _02107_ reset_n keymem.key_mem\[0\]\[71\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22826_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[125\] _06839_ _03864_ _05085_ _02161_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_211_1410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25545_ VGND VPWR VPWR VGND clk _02038_ reset_n keymem.key_mem\[0\]\[2\] sky130_fd_sc_hd__dfrtp_2
X_22757_ VGND VPWR _02109_ _06843_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12510_ VGND VPWR _08077_ _07551_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_26_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13490_ VPWR VGND VPWR VGND _08962_ enc_block.block_w0_reg\[3\] _08952_ sky130_fd_sc_hd__or2_2
X_21708_ VGND VPWR _01580_ _06323_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25476_ VGND VPWR VPWR VGND clk _01969_ reset_n keymem.key_mem\[1\]\[61\] sky130_fd_sc_hd__dfrtp_2
X_22688_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[32\] _06790_ _06789_ _04920_ _02068_
+ sky130_fd_sc_hd__a22o_2
X_12441_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[29\] _07893_ _08014_ _08007_ _08015_
+ sky130_fd_sc_hd__o22a_2
X_24427_ VGND VPWR VPWR VGND clk _00920_ reset_n keymem.key_mem\[9\]\[36\] sky130_fd_sc_hd__dfrtp_2
X_21639_ VGND VPWR _01547_ _06287_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_30_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15160_ VPWR VGND VGND VPWR _10562_ _10623_ _10611_ _10624_ sky130_fd_sc_hd__nor3_2
XFILLER_0_34_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12372_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[23\] _07535_ _07951_ _07945_ _07952_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_129_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24358_ VGND VPWR VPWR VGND clk _00851_ reset_n keymem.key_mem\[10\]\[95\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_164_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14111_ VGND VPWR _09582_ _09340_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_65_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15091_ VGND VPWR VGND VPWR _10520_ _10554_ _10469_ _10475_ _10553_ _10555_ sky130_fd_sc_hd__o32a_2
XFILLER_0_26_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23309_ VGND VPWR VGND VPWR _07189_ _04505_ _07187_ _07188_ _07190_ sky130_fd_sc_hd__a31o_2
XPHY_EDGE_ROW_135_1_Right_736 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24289_ VGND VPWR VPWR VGND clk _00782_ reset_n keymem.key_mem\[10\]\[26\] sky130_fd_sc_hd__dfrtp_2
X_14042_ VGND VPWR _09514_ _09513_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18850_ VGND VPWR VGND VPWR _04694_ _04693_ _04696_ _04692_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_66_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17801_ VGND VPWR VGND VPWR _03134_ _03792_ _03795_ _03793_ _03727_ _03797_ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_98_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18781_ VPWR VGND VGND VPWR _04613_ _04634_ _04019_ sky130_fd_sc_hd__nor2_2
X_15993_ VGND VPWR _00028_ _11448_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_179_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_101_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17732_ VGND VPWR VPWR VGND _03723_ _02880_ keymem.prev_key0_reg\[33\] _03754_ sky130_fd_sc_hd__mux2_2
X_14944_ VGND VPWR VGND VPWR _10408_ _10407_ _10406_ keymem.prev_key1_reg\[11\] _08955_
+ _08942_ sky130_fd_sc_hd__a32o_2
XFILLER_0_76_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_89_315 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_136_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17663_ VGND VPWR VPWR VGND _03691_ key[141] keymem.prev_key1_reg\[13\] _03705_ sky130_fd_sc_hd__mux2_2
X_14875_ VGND VPWR VPWR VGND _09036_ _09129_ _09041_ _10340_ sky130_fd_sc_hd__or3_2
XFILLER_0_72_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_833 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_76_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19402_ VPWR VGND keymem.key_mem\[12\]\[1\] _05097_ _05095_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_159_214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16614_ VGND VPWR VPWR VGND _02769_ _02770_ _07387_ _02767_ _02768_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_159_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13826_ VGND VPWR VGND VPWR _09298_ _09259_ _09258_ keymem.prev_key1_reg\[26\] _08989_
+ _08983_ sky130_fd_sc_hd__a32o_2
XFILLER_0_106_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17594_ VPWR VGND VPWR VGND _03651_ _10323_ _03653_ _03652_ keylen sky130_fd_sc_hd__a211oi_2
X_19333_ VGND VPWR _00479_ _05049_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16545_ VGND VPWR _02704_ keymem.prev_key0_reg\[25\] _02703_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_13757_ VPWR VGND VGND VPWR _09228_ _09108_ _09229_ _09082_ _09095_ _09157_ sky130_fd_sc_hd__o32ai_2
XFILLER_0_202_398 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_57_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_919 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_174_228 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12708_ VGND VPWR VGND VPWR _08096_ keymem.key_mem\[5\]\[54\] _08253_ _08255_ _08257_
+ _08256_ sky130_fd_sc_hd__a2111o_2
X_19264_ VPWR VGND keymem.key_mem\[13\]\[83\] _05005_ _04979_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16476_ VPWR VGND VGND VPWR _02613_ _02620_ _02636_ _02637_ sky130_fd_sc_hd__nor3_2
X_13688_ VGND VPWR _09160_ _09159_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_57_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18215_ VPWR VGND _04124_ _04123_ enc_block.round_key\[109\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15427_ VPWR VGND VGND VPWR _10535_ _10574_ _10888_ _10575_ _10635_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_122_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12639_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[48\] _07744_ keymem.key_mem\[10\]\[48\]
+ _08193_ _08194_ sky130_fd_sc_hd__a22o_2
X_19195_ VGND VPWR VPWR VGND _04951_ _04963_ keymem.key_mem\[13\]\[55\] _04964_ sky130_fd_sc_hd__mux2_2
XFILLER_0_26_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_963 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_127_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_147_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_186_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18146_ VPWR VGND _04061_ _04060_ enc_block.round_key\[103\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_83_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_53_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15358_ VGND VPWR VGND VPWR _10818_ _10817_ _10820_ _10819_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_14_838 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_87_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_147_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14309_ VPWR VGND VPWR VGND _09772_ _09778_ _09775_ _09771_ _09779_ sky130_fd_sc_hd__or4_2
XFILLER_0_83_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18077_ VPWR VGND _03997_ enc_block.block_w0_reg\[25\] enc_block.block_w3_reg\[1\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_44_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15289_ VGND VPWR _10751_ _10557_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_1_732 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_262_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17028_ VGND VPWR _00072_ _03151_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_106_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_226_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_77_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18979_ VPWR VGND VPWR VGND _04811_ block[55] _04744_ enc_block.block_w3_reg\[23\]
+ _04798_ _04812_ sky130_fd_sc_hd__a221o_2
XFILLER_0_225_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_457 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_193_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21990_ VGND VPWR _06475_ _06403_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_94_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_154_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20941_ VGND VPWR VGND VPWR _05917_ keymem.key_mem_we _03322_ _05916_ _01219_ sky130_fd_sc_hd__a31o_2
XFILLER_0_193_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20872_ VGND VPWR _05880_ _05819_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_221_663 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23660_ keymem.prev_key0_reg\[16\] clk _00157_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_7_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22611_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[121\] _06777_ _06776_ _05077_ _02029_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_7_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_810 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23591_ VGND VPWR VPWR VGND clk _00092_ reset_n keymem.key_mem\[14\]\[80\] sky130_fd_sc_hd__dfrtp_2
X_22542_ VGND VPWR VPWR VGND _06750_ keymem.key_mem\[1\]\[71\] _03252_ _06759_ sky130_fd_sc_hd__mux2_2
X_25330_ VGND VPWR VPWR VGND clk _01823_ reset_n keymem.key_mem\[2\]\[43\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_178_2_Right_250 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_130_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22473_ VGND VPWR VPWR VGND _06726_ keymem.key_mem\[1\]\[30\] _02839_ _06731_ sky130_fd_sc_hd__mux2_2
X_25261_ VGND VPWR VPWR VGND clk _01754_ reset_n keymem.key_mem\[3\]\[102\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_165_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21424_ VGND VPWR _06173_ _06116_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24212_ VGND VPWR VPWR VGND clk _00705_ reset_n keymem.key_mem\[11\]\[77\] sky130_fd_sc_hd__dfrtp_2
X_25192_ VGND VPWR VPWR VGND clk _01685_ reset_n keymem.key_mem\[3\]\[33\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_165_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_245_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24143_ VGND VPWR VPWR VGND clk _00636_ reset_n keymem.key_mem\[11\]\[8\] sky130_fd_sc_hd__dfrtp_2
X_21355_ VGND VPWR VPWR VGND _06128_ _02339_ keymem.key_mem\[5\]\[18\] _06137_ sky130_fd_sc_hd__mux2_2
XFILLER_0_62_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_114_394 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20306_ VGND VPWR _00923_ _05578_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24074_ VGND VPWR VPWR VGND clk _00567_ reset_n keymem.key_mem\[12\]\[67\] sky130_fd_sc_hd__dfrtp_2
X_21286_ VGND VPWR _01382_ _06099_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_13_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_241_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_690 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23025_ VPWR VGND VPWR VGND _06982_ keymem.prev_key1_reg\[62\] _06926_ sky130_fd_sc_hd__or2_2
X_20237_ VGND VPWR _00890_ _05542_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_229_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_102_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20168_ VGND VPWR _05504_ _05387_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12990_ VGND VPWR VGND VPWR _08511_ _07690_ keymem.key_mem\[3\]\[82\] _08510_ _07746_
+ sky130_fd_sc_hd__a211o_2
X_20099_ VGND VPWR VPWR VGND _05457_ _03252_ keymem.key_mem\[10\]\[71\] _05468_ sky130_fd_sc_hd__mux2_2
X_24976_ VGND VPWR VPWR VGND clk _01469_ reset_n keymem.key_mem\[5\]\[73\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_172_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23927_ VGND VPWR VPWR VGND clk _00420_ reset_n keymem.key_mem\[13\]\[48\] sky130_fd_sc_hd__dfrtp_2
X_11941_ VPWR VGND VGND VPWR _07543_ _07544_ _07530_ sky130_fd_sc_hd__nor2_2
XFILLER_0_19_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_231_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_197_821 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_213_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14660_ VPWR VGND VPWR VGND _10045_ _10126_ _10123_ _09899_ _10127_ sky130_fd_sc_hd__or4_2
XFILLER_0_54_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23858_ VGND VPWR VPWR VGND clk _00351_ reset_n enc_block.block_w2_reg\[11\] sky130_fd_sc_hd__dfrtp_2
X_11872_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[7\] dec_new_block\[103\]
+ _07500_ sky130_fd_sc_hd__mux2_2
XFILLER_0_211_140 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_197_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13611_ VGND VPWR VGND VPWR _09083_ _09039_ _09041_ _09057_ _09010_ sky130_fd_sc_hd__a211o_2
XFILLER_0_213_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_696 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22809_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[110\] _06858_ _06857_ _05054_ _02146_
+ sky130_fd_sc_hd__a22o_2
X_14591_ VPWR VGND VPWR VGND _10057_ _10058_ _10059_ _09579_ _09911_ sky130_fd_sc_hd__or4b_2
X_23789_ VGND VPWR VPWR VGND clk _00282_ reset_n enc_block.block_w0_reg\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_200_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16330_ VGND VPWR VPWR VGND _02493_ keymem.prev_key1_reg\[53\] _02491_ _02492_ _08927_
+ sky130_fd_sc_hd__o31a_2
X_13542_ VGND VPWR _09014_ _09013_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25528_ VGND VPWR VPWR VGND clk _02021_ reset_n keymem.key_mem\[1\]\[113\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_429 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16261_ VPWR VGND VPWR VGND _02424_ _11503_ _11365_ _11596_ _11417_ _02425_ sky130_fd_sc_hd__a221o_2
XFILLER_0_54_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13473_ VGND VPWR _08945_ _08944_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25459_ VGND VPWR VPWR VGND clk _01952_ reset_n keymem.key_mem\[1\]\[44\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_246_1325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18000_ VPWR VGND VPWR VGND _03932_ _03729_ _03931_ sky130_fd_sc_hd__or2_2
X_15212_ VGND VPWR VPWR VGND _10516_ _10545_ _10515_ _10675_ sky130_fd_sc_hd__or3_2
X_12424_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[28\] _07602_ keymem.key_mem\[7\]\[28\]
+ _07567_ _07999_ sky130_fd_sc_hd__a22o_2
X_16192_ VGND VPWR VGND VPWR _11308_ _11465_ _11204_ _11385_ _02357_ sky130_fd_sc_hd__o22a_2
XFILLER_0_129_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_50_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_69_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15143_ VGND VPWR VGND VPWR _10521_ _10566_ _10513_ _10593_ _10607_ sky130_fd_sc_hd__o22a_2
XFILLER_0_51_966 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_105_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12355_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[22\] _07586_ keymem.key_mem\[6\]\[22\]
+ _07564_ _07936_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_136_1_Right_737 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15074_ VGND VPWR _10538_ _10484_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12286_ VGND VPWR _07872_ _07567_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19951_ VGND VPWR _00756_ _05390_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_220_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_2_Left_575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_267_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14025_ VPWR VGND VGND VPWR _09496_ _09493_ _09447_ _09360_ _09464_ _09497_ sky130_fd_sc_hd__a311o_2
X_18902_ VPWR VGND VGND VPWR _04654_ _04743_ _04137_ sky130_fd_sc_hd__nor2_2
XFILLER_0_120_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19882_ VGND VPWR _00725_ _05352_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_208_914 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_208_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_73_1_Left_340 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18833_ VGND VPWR VGND VPWR _04679_ enc_block.round_key\[40\] _04681_ _04266_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_184_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_93_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18764_ VPWR VGND VPWR VGND _04618_ _04615_ _04617_ sky130_fd_sc_hd__or2_2
XFILLER_0_218_1416 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15976_ VGND VPWR VGND VPWR _11432_ _11229_ _11289_ _11272_ _11288_ sky130_fd_sc_hd__and4_2
X_17715_ VGND VPWR VGND VPWR _03732_ keymem.prev_key1_reg\[27\] _03743_ _03733_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_37_1202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14927_ VPWR VGND VPWR VGND _10391_ enc_block.block_w0_reg\[9\] _09273_ sky130_fd_sc_hd__or2_2
XFILLER_0_76_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18695_ _04554_ _04556_ _04294_ _04555_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_26_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17646_ VGND VPWR _00148_ _03693_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_158_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14858_ VGND VPWR _10323_ _10322_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_118_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13809_ enc_block.sword_ctr_reg\[1\] _09281_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[29\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_216_1195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_4_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1086 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17577_ VPWR VGND VGND VPWR _11456_ _03638_ key[251] sky130_fd_sc_hd__nor2_2
X_14789_ VGND VPWR VGND VPWR _10255_ _10254_ _10253_ _10252_ _10251_ sky130_fd_sc_hd__and4_2
X_19316_ VGND VPWR VPWR VGND _05025_ _05037_ keymem.key_mem\[13\]\[102\] _05038_ sky130_fd_sc_hd__mux2_2
XFILLER_0_42_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16528_ VPWR VGND VPWR VGND _02687_ _02677_ _02676_ key[152] _11043_ _02688_ sky130_fd_sc_hd__a221o_2
XFILLER_0_45_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_42_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19247_ VGND VPWR _00448_ _04994_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16459_ VPWR VGND VPWR VGND _02616_ _02619_ _02617_ _11431_ _02620_ sky130_fd_sc_hd__or4_2
XFILLER_0_186_1261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_42_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19178_ VPWR VGND keymem.key_mem_we _04953_ _03046_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_83_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_87_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18129_ VGND VPWR _04045_ enc_block.block_w3_reg\[5\] enc_block.block_w0_reg\[29\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_147_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_83_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_48_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21140_ VGND VPWR VPWR VGND _06018_ _03006_ keymem.key_mem\[6\]\[45\] _06023_ sky130_fd_sc_hd__mux2_2
XFILLER_0_223_1133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_258_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_223_1177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_158_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21071_ VGND VPWR VPWR VGND _05983_ _10976_ keymem.key_mem\[6\]\[12\] _05987_ sky130_fd_sc_hd__mux2_2
XFILLER_0_10_874 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20022_ VGND VPWR VPWR VGND _05424_ _02894_ keymem.key_mem\[10\]\[34\] _05428_ sky130_fd_sc_hd__mux2_2
XFILLER_0_158_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24830_ VGND VPWR VPWR VGND clk _01323_ reset_n keymem.key_mem\[6\]\[55\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_158_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24761_ VGND VPWR VPWR VGND clk _01254_ reset_n keymem.key_mem\[7\]\[114\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_154_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21973_ VPWR VGND keymem.key_mem\[3\]\[51\] _06466_ _06439_ VPWR VGND sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_61_Left_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_59_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23712_ keymem.prev_key0_reg\[68\] clk _00209_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_94_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20924_ VGND VPWR VPWR VGND _05880_ _04986_ keymem.key_mem\[7\]\[72\] _05908_ sky130_fd_sc_hd__mux2_2
XFILLER_0_55_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24692_ VGND VPWR VPWR VGND clk _01185_ reset_n keymem.key_mem\[7\]\[45\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_7_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20855_ VGND VPWR _01179_ _05871_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23643_ VGND VPWR VPWR VGND clk _00003_ reset_n keymem.ready_new sky130_fd_sc_hd__dfrtp_2
XFILLER_0_193_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23574_ VGND VPWR VPWR VGND clk _00075_ reset_n keymem.key_mem\[14\]\[63\] sky130_fd_sc_hd__dfrtp_2
X_20786_ VPWR VGND keymem.key_mem\[7\]\[8\] _05834_ _05830_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_153_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25313_ VGND VPWR VPWR VGND clk _01806_ reset_n keymem.key_mem\[2\]\[26\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_64_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22525_ VGND VPWR _06750_ _06695_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_179_2_Right_251 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_106_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25244_ VGND VPWR VPWR VGND clk _01737_ reset_n keymem.key_mem\[3\]\[85\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_165_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22456_ VGND VPWR VPWR VGND _06715_ keymem.key_mem\[1\]\[22\] _02608_ _06722_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_484 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_32_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_66_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21407_ VGND VPWR _01438_ _06164_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25175_ VGND VPWR VPWR VGND clk _01668_ reset_n keymem.key_mem\[3\]\[16\] sky130_fd_sc_hd__dfrtp_2
X_22387_ VGND VPWR VPWR VGND _06680_ _03607_ keymem.key_mem\[2\]\[118\] _06685_ sky130_fd_sc_hd__mux2_2
XFILLER_0_66_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12140_ VPWR VGND VPWR VGND _07735_ keymem.key_mem\[13\]\[7\] _07731_ keymem.key_mem\[3\]\[7\]
+ _07691_ _07736_ sky130_fd_sc_hd__a221o_2
X_24126_ VGND VPWR VPWR VGND clk _00619_ reset_n keymem.key_mem\[12\]\[119\] sky130_fd_sc_hd__dfrtp_2
X_21338_ VGND VPWR _06128_ _06116_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_13_690 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1277 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12071_ VGND VPWR _07671_ _07670_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24057_ VGND VPWR VPWR VGND clk _00550_ reset_n keymem.key_mem\[12\]\[50\] sky130_fd_sc_hd__dfrtp_2
X_21269_ VGND VPWR _01374_ _06090_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1143 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_263_316 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23008_ VGND VPWR VGND VPWR _03094_ _03093_ _03098_ _06972_ sky130_fd_sc_hd__a21o_2
XFILLER_0_102_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15830_ VGND VPWR _11286_ _11247_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_102_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_265 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_176_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_736 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15761_ VPWR VGND VPWR VGND _11172_ _11216_ _11179_ _11166_ _11217_ sky130_fd_sc_hd__or4_2
XFILLER_0_77_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24959_ VGND VPWR VPWR VGND clk _01452_ reset_n keymem.key_mem\[5\]\[56\] sky130_fd_sc_hd__dfrtp_2
X_12973_ VGND VPWR enc_block.round_key\[80\] _08495_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_137_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17500_ VGND VPWR VPWR VGND _09927_ _11452_ key[241] _03571_ sky130_fd_sc_hd__mux2_2
X_14712_ VPWR VGND VGND VPWR _09141_ _10179_ _09153_ sky130_fd_sc_hd__nor2_2
XFILLER_0_73_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18480_ VGND VPWR _04363_ enc_block.block_w3_reg\[13\] enc_block.block_w2_reg\[21\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_11924_ VPWR VGND VPWR VGND _07527_ _07525_ _07526_ sky130_fd_sc_hd__or2_2
X_15692_ VGND VPWR _11149_ _11148_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_217_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_611 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_234_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17431_ VGND VPWR VPWR VGND _03467_ keymem.key_mem\[14\]\[103\] _03511_ _03512_ sky130_fd_sc_hd__mux2_2
XFILLER_0_197_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14643_ VPWR VGND VPWR VGND _09599_ _09603_ _10109_ _09432_ _10110_ sky130_fd_sc_hd__or4_2
X_11855_ VGND VPWR result[94] _07491_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_86_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_135_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_196_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_513 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17362_ VPWR VGND VPWR VGND _03451_ _10902_ _03449_ key[222] _03366_ _03452_ sky130_fd_sc_hd__a221o_2
X_14574_ VGND VPWR VGND VPWR _09327_ _09415_ _09305_ _09411_ _10042_ sky130_fd_sc_hd__o22a_2
XFILLER_0_71_1192 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11786_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[28\] dec_new_block\[60\]
+ _07457_ sky130_fd_sc_hd__mux2_2
XFILLER_0_32_1154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19101_ VGND VPWR VGND VPWR _04905_ keymem.key_mem_we _02410_ _04896_ _00391_ sky130_fd_sc_hd__a31o_2
XFILLER_0_144_209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16313_ VPWR VGND VGND VPWR _02476_ _02477_ _02475_ sky130_fd_sc_hd__nor2_2
X_13525_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[4\] _08969_ _08997_ _08964_ _08994_
+ _08996_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_113_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17293_ VPWR VGND VPWR VGND _03390_ key[87] _09795_ sky130_fd_sc_hd__or2_2
XFILLER_0_250_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19032_ VGND VPWR _04859_ enc_block.round_key\[61\] _04858_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16244_ VPWR VGND VPWR VGND _02408_ _02401_ _02343_ key[147] _11043_ _02409_ sky130_fd_sc_hd__a221o_2
XFILLER_0_183_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13456_ VPWR VGND VGND VPWR _08927_ _08928_ _07378_ sky130_fd_sc_hd__nor2_2
XFILLER_0_148_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_144_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12407_ VGND VPWR enc_block.round_key\[26\] _07983_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_88_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16175_ VGND VPWR VPWR VGND _11041_ keymem.key_mem\[14\]\[18\] _02340_ _02341_ sky130_fd_sc_hd__mux2_2
X_13387_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[122\] _07659_ keymem.key_mem\[7\]\[122\]
+ _07608_ _08868_ sky130_fd_sc_hd__a22o_2
XFILLER_0_2_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15126_ VPWR VGND VGND VPWR _10500_ _10590_ _10472_ sky130_fd_sc_hd__nor2_2
XFILLER_0_45_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_224_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12338_ VGND VPWR VGND VPWR _07921_ _07919_ keymem.key_mem\[9\]\[20\] _07920_ _07572_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_266_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_137_1_Right_738 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15057_ VGND VPWR _10521_ _10414_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_259_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_267_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19934_ VGND VPWR _00750_ _05379_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12269_ VPWR VGND VPWR VGND _07856_ keymem.key_mem\[9\]\[15\] _07672_ keymem.key_mem\[4\]\[15\]
+ _07854_ _07857_ sky130_fd_sc_hd__a221o_2
X_14008_ VGND VPWR _09480_ _09329_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_259_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19865_ VGND VPWR _00717_ _05343_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_120_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18816_ VPWR VGND VPWR VGND _04665_ _04664_ _04663_ enc_block.block_w2_reg\[6\] _04602_
+ _00346_ sky130_fd_sc_hd__a221o_2
X_19796_ VGND VPWR _00684_ _05307_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_155_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_222_Left_489 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_194_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15959_ VPWR VGND VPWR VGND _11411_ _11414_ _11413_ _11410_ _11415_ sky130_fd_sc_hd__or4_2
X_18747_ VGND VPWR _04602_ _04599_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_222_224 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_155_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18678_ VPWR VGND _04541_ _04540_ enc_block.round_key\[89\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_77_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_231_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1065 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_8_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17629_ VGND VPWR VPWR VGND _03681_ _03680_ keymem.prev_key0_reg\[2\] _03682_ sky130_fd_sc_hd__mux2_2
XFILLER_0_231_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_323 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20640_ VGND VPWR _01081_ _05754_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_175_345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_1254 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_266_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_343 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20571_ VGND VPWR _01048_ _05718_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_188_1389 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22310_ VGND VPWR _01861_ _06644_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_231_Left_498 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23290_ VPWR VGND _07173_ _07172_ enc_block.round_key\[8\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_61_527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_1085 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_944 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_14_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_1_Right_700 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_82_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22241_ VGND VPWR _01828_ _06608_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_162_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1228 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_15_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22172_ VGND VPWR _01795_ _06572_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_169_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_242_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21123_ VGND VPWR VPWR VGND _06007_ _02923_ keymem.key_mem\[6\]\[37\] _06014_ sky130_fd_sc_hd__mux2_2
XFILLER_0_203_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_143 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_218_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_95 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_160_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21054_ VGND VPWR _01272_ _05977_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_258_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20005_ VGND VPWR VPWR VGND _05413_ _02743_ keymem.key_mem\[10\]\[26\] _05419_ sky130_fd_sc_hd__mux2_2
XFILLER_0_226_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_94_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24813_ VGND VPWR VPWR VGND clk _01306_ reset_n keymem.key_mem\[6\]\[38\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_158_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25793_ keymem.prev_key1_reg\[109\] clk _02286_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_55_1121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24744_ VGND VPWR VPWR VGND clk _01237_ reset_n keymem.key_mem\[7\]\[97\] sky130_fd_sc_hd__dfrtp_2
X_21956_ VGND VPWR VPWR VGND _06449_ _04941_ keymem.key_mem\[3\]\[43\] _06457_ sky130_fd_sc_hd__mux2_2
XFILLER_0_201_419 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20907_ VGND VPWR _05899_ _05822_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_178_161 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24675_ VGND VPWR VPWR VGND clk _01168_ reset_n keymem.key_mem\[7\]\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21887_ VGND VPWR _01663_ _06419_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23626_ VGND VPWR VPWR VGND clk _00127_ reset_n keymem.key_mem\[14\]\[115\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_166_345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11640_ VGND VPWR VGND VPWR enc_block.round\[1\] enc_block.round\[2\] _07378_ _07379_
+ sky130_fd_sc_hd__a21o_2
X_20838_ VGND VPWR VPWR VGND _05820_ _04920_ keymem.key_mem\[7\]\[32\] _05862_ sky130_fd_sc_hd__mux2_2
XFILLER_0_64_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_119_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23557_ VGND VPWR VPWR VGND clk _00058_ reset_n keymem.key_mem\[14\]\[46\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_64_354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20769_ VPWR VGND keymem.key_mem\[7\]\[0\] _05825_ _05824_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_181_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_64_376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_294 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13310_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[114\] _07924_ keymem.key_mem\[10\]\[114\]
+ _07876_ _08799_ sky130_fd_sc_hd__a22o_2
XFILLER_0_24_218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22508_ VGND VPWR VPWR VGND _06739_ keymem.key_mem\[1\]\[54\] _03091_ _06742_ sky130_fd_sc_hd__mux2_2
X_14290_ VPWR VGND VGND VPWR _09348_ _09403_ _09760_ _09311_ _09563_ sky130_fd_sc_hd__o22ai_2
X_23488_ VPWR VGND VPWR VGND _07349_ _03950_ _07348_ enc_block.block_w3_reg\[29\]
+ _07126_ _02334_ sky130_fd_sc_hd__a221o_2
XFILLER_0_134_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_257_Right_126 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25227_ VGND VPWR VPWR VGND clk _01720_ reset_n keymem.key_mem\[3\]\[68\] sky130_fd_sc_hd__dfrtp_2
X_13241_ VGND VPWR VGND VPWR _07786_ keymem.key_mem\[10\]\[107\] _08733_ _08735_ _08737_
+ _08736_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_21_903 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22439_ VGND VPWR VPWR VGND _06702_ keymem.key_mem\[1\]\[14\] _11099_ _06713_ sky130_fd_sc_hd__mux2_2
XFILLER_0_27_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_66_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13172_ VGND VPWR VGND VPWR _08675_ _07588_ keymem.key_mem\[13\]\[100\] _08674_ _07616_
+ sky130_fd_sc_hd__a211o_2
X_25158_ VGND VPWR VPWR VGND clk _01651_ reset_n keymem.key_mem\[4\]\[127\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24109_ VGND VPWR VPWR VGND clk _00602_ reset_n keymem.key_mem\[12\]\[102\] sky130_fd_sc_hd__dfrtp_2
X_12123_ VGND VPWR VGND VPWR _07712_ keymem.key_mem\[6\]\[6\] _07713_ _07719_ _07720_
+ _07663_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_27_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17980_ VGND VPWR _00257_ _03918_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_20_468 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25089_ VGND VPWR VPWR VGND clk _01582_ reset_n keymem.key_mem\[4\]\[58\] sky130_fd_sc_hd__dfrtp_2
X_16931_ VPWR VGND VPWR VGND _03064_ keymem.prev_key1_reg\[51\] sky130_fd_sc_hd__inv_2
XFILLER_0_263_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12054_ VGND VPWR _07654_ _07538_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_245_850 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16862_ VGND VPWR VGND VPWR _03001_ _02928_ _02927_ key[45] sky130_fd_sc_hd__o21a_2
X_19650_ VGND VPWR VPWR VGND _05227_ _05069_ keymem.key_mem\[12\]\[117\] _05229_ sky130_fd_sc_hd__mux2_2
XFILLER_0_74_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15813_ VGND VPWR VPWR VGND _11265_ _11180_ _11167_ _11269_ sky130_fd_sc_hd__or3_2
X_18601_ VGND VPWR _04472_ _04401_ _04471_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_254_1424 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_137_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19581_ VGND VPWR VPWR VGND _05183_ _05006_ keymem.key_mem\[12\]\[84\] _05193_ sky130_fd_sc_hd__mux2_2
X_16793_ VGND VPWR VGND VPWR _02938_ _09512_ _11543_ key[39] sky130_fd_sc_hd__o21a_2
XFILLER_0_99_251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18532_ VGND VPWR _04410_ enc_block.block_w3_reg\[9\] enc_block.block_w1_reg\[26\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_232_566 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_137_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15744_ VGND VPWR VGND VPWR enc_block.block_w1_reg\[21\] _08985_ _10387_ _11198_
+ _11200_ _11199_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_38_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12956_ VGND VPWR _08480_ _07746_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_34_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11907_ VGND VPWR result[120] _07517_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18463_ VGND VPWR VGND VPWR _04347_ _04065_ _04345_ _04346_ _04348_ sky130_fd_sc_hd__a31o_2
XFILLER_0_59_148 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_213_791 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15675_ VGND VPWR VGND VPWR _10667_ _10751_ _10482_ _10867_ _11132_ sky130_fd_sc_hd__o22a_2
XFILLER_0_114_13 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12887_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[72\] _07609_ keymem.key_mem\[8\]\[72\]
+ _07929_ _08418_ sky130_fd_sc_hd__a22o_2
XFILLER_0_213_1154 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17414_ VGND VPWR VPWR VGND _09732_ _10142_ key[229] _03497_ sky130_fd_sc_hd__mux2_2
X_14626_ VGND VPWR VGND VPWR _10094_ _10093_ _10090_ _09522_ sky130_fd_sc_hd__o21a_2
X_11838_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[22\] dec_new_block\[86\]
+ _07483_ sky130_fd_sc_hd__mux2_2
X_18394_ VPWR VGND VPWR VGND _04286_ _04044_ _04285_ sky130_fd_sc_hd__or2_2
XFILLER_0_67_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_153 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17345_ VGND VPWR _00104_ _03436_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_184_175 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_150_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14557_ VPWR VGND VGND VPWR _09153_ _10025_ _09090_ sky130_fd_sc_hd__nor2_2
X_11769_ VGND VPWR result[51] _07448_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_28_579 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_43_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_82_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13508_ VPWR VGND VPWR VGND _08979_ _08948_ _08978_ _08945_ enc_block.block_w2_reg\[6\]
+ _08980_ sky130_fd_sc_hd__a221o_2
X_17276_ VGND VPWR VPWR VGND _03296_ keymem.key_mem\[14\]\[85\] _03374_ _03375_ sky130_fd_sc_hd__mux2_2
X_14488_ VPWR VGND VGND VPWR _09077_ _09112_ _09957_ _09134_ _09036_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_3_602 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_148_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19015_ VPWR VGND _04844_ _04843_ enc_block.round_key\[59\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_183_1242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16227_ VPWR VGND VPWR VGND _02388_ _02391_ _02392_ _02384_ _11322_ sky130_fd_sc_hd__or4b_2
X_13439_ VGND VPWR VGND VPWR _07780_ keymem.key_mem\[5\]\[127\] _08912_ _08914_ _08915_
+ _07573_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_109_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_796 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16158_ VPWR VGND VGND VPWR _11403_ _11612_ _11298_ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_947 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15109_ VPWR VGND VPWR VGND _10473_ _10466_ _10440_ _10451_ _10573_ sky130_fd_sc_hd__or4_2
XFILLER_0_239_143 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16089_ VPWR VGND VPWR VGND _11544_ key[17] _11543_ sky130_fd_sc_hd__or2_2
XFILLER_0_48_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_1_Right_739 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19917_ VGND VPWR _00742_ _05370_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_48_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_259_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19848_ VGND VPWR _00709_ _05334_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_39_1116 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_194_1360 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_155_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19779_ VGND VPWR _00676_ _05298_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_190_1213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_223_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21810_ VGND VPWR _01629_ _06376_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_56_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22790_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[94\] _06850_ _06849_ _05021_ _02130_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_210_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_116_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21741_ VGND VPWR _01596_ _06340_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_8_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_811 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_129_2_Left_600 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24460_ VGND VPWR VPWR VGND clk _00953_ reset_n keymem.key_mem\[9\]\[69\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_524 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21672_ VGND VPWR _01563_ _06304_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_46_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23411_ VPWR VGND VGND VPWR _07192_ _07282_ _04201_ sky130_fd_sc_hd__nor2_2
XFILLER_0_266_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20623_ VGND VPWR _01073_ _05745_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_163_326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24391_ VGND VPWR VPWR VGND clk _00884_ reset_n keymem.key_mem\[9\]\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_163_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1057 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23342_ VGND VPWR VGND VPWR _07219_ _03949_ _04125_ _07220_ sky130_fd_sc_hd__a21o_2
X_20554_ VGND VPWR _01040_ _05709_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_116_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_62_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_166_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23273_ VGND VPWR _07157_ enc_block.block_w3_reg\[31\] enc_block.block_w0_reg\[23\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20485_ VGND VPWR VPWR VGND _05534_ _03654_ keymem.key_mem\[9\]\[125\] _05672_ sky130_fd_sc_hd__mux2_2
XFILLER_0_63_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25012_ VGND VPWR VPWR VGND clk _01505_ reset_n keymem.key_mem\[5\]\[109\] sky130_fd_sc_hd__dfrtp_2
X_22224_ VGND VPWR _01820_ _06599_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_28_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22155_ VGND VPWR VPWR VGND _06554_ _10661_ keymem.key_mem\[2\]\[8\] _06563_ sky130_fd_sc_hd__mux2_2
XFILLER_0_24_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21106_ VGND VPWR VPWR VGND _05996_ _02811_ keymem.key_mem\[6\]\[29\] _06005_ sky130_fd_sc_hd__mux2_2
XFILLER_0_98_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22086_ VGND VPWR _01756_ _06525_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_238_1419 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21037_ VGND VPWR VPWR VGND _05819_ _05087_ keymem.key_mem\[7\]\[126\] _05967_ sky130_fd_sc_hd__mux2_2
XFILLER_0_261_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_22_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_138_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_864 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12810_ VGND VPWR VGND VPWR _08349_ _07968_ keymem.key_mem\[9\]\[64\] _08346_ _08348_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_242_886 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1007 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13790_ VGND VPWR VGND VPWR _09262_ enc_block.block_w2_reg\[25\] enc_block.sword_ctr_reg\[1\]
+ enc_block.sword_ctr_reg\[0\] sky130_fd_sc_hd__and3b_2
X_25776_ keymem.prev_key1_reg\[92\] clk _02269_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22988_ VGND VPWR VPWR VGND _06960_ _06959_ keymem.prev_key1_reg\[46\] _06961_ sky130_fd_sc_hd__mux2_2
XFILLER_0_74_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24727_ VGND VPWR VPWR VGND clk _01220_ reset_n keymem.key_mem\[7\]\[80\] sky130_fd_sc_hd__dfrtp_2
X_12741_ VGND VPWR VGND VPWR _07793_ keymem.key_mem\[0\]\[57\] _08286_ _08281_ _08279_
+ _08287_ sky130_fd_sc_hd__o32a_2
XFILLER_0_214_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21939_ VPWR VGND keymem.key_mem\[3\]\[35\] _06448_ _06439_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_139_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_750 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15460_ VPWR VGND VPWR VGND _10752_ _10919_ _10777_ _10918_ _10920_ sky130_fd_sc_hd__or4_2
XFILLER_0_214_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12672_ VPWR VGND VPWR VGND _08223_ keymem.key_mem\[6\]\[51\] _07739_ keymem.key_mem\[10\]\[51\]
+ _07865_ _08224_ sky130_fd_sc_hd__a221o_2
X_24658_ VGND VPWR VPWR VGND clk _01151_ reset_n keymem.key_mem\[7\]\[11\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_113_2_Left_584 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14411_ VPWR VGND VGND VPWR _09353_ _09381_ _09880_ _09389_ _09415_ sky130_fd_sc_hd__o22ai_2
X_23609_ VGND VPWR VPWR VGND clk _00110_ reset_n keymem.key_mem\[14\]\[98\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_249_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15391_ VPWR VGND VGND VPWR _10644_ _10852_ _10595_ sky130_fd_sc_hd__nor2_2
XFILLER_0_37_354 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24589_ VGND VPWR VPWR VGND clk _01082_ reset_n keymem.key_mem\[8\]\[70\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_166_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17130_ VGND VPWR VGND VPWR _03243_ _10277_ _03244_ keylen sky130_fd_sc_hd__a21oi_2
X_14342_ VGND VPWR VGND VPWR _09812_ _09153_ _09110_ _09687_ _09211_ _09811_ sky130_fd_sc_hd__o221ai_2
X_17061_ VPWR VGND VPWR VGND _03182_ _10086_ _03179_ _03180_ _03181_ _10096_ sky130_fd_sc_hd__o311a_2
XFILLER_0_162_370 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14273_ VGND VPWR VPWR VGND _09339_ _09309_ _09306_ _09743_ sky130_fd_sc_hd__or3_2
XFILLER_0_145_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16012_ VPWR VGND VGND VPWR _11380_ _11379_ _11467_ _11466_ _11464_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_21_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13224_ VGND VPWR VGND VPWR _08722_ _07808_ keymem.key_mem\[12\]\[105\] _08719_ _08721_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_106_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_278 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13155_ VGND VPWR enc_block.round_key\[98\] _08659_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12106_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[5\] _07597_ keymem.key_mem\[7\]\[5\]
+ _07703_ _07704_ sky130_fd_sc_hd__a22o_2
X_17963_ VGND VPWR VPWR VGND _03896_ _03906_ keymem.prev_key0_reg\[111\] _03907_ sky130_fd_sc_hd__mux2_2
X_13086_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[92\] _07872_ keymem.key_mem\[2\]\[92\]
+ _07697_ _08597_ sky130_fd_sc_hd__a22o_2
XFILLER_0_256_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19702_ VGND VPWR VPWR VGND _05247_ keymem.key_mem\[11\]\[12\] _10977_ _05258_ sky130_fd_sc_hd__mux2_2
X_16914_ VPWR VGND VGND VPWR _02947_ _11560_ _11622_ _03048_ sky130_fd_sc_hd__nor3_2
X_12037_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[2\] _07603_ keymem.key_mem\[4\]\[2\]
+ _07637_ _07638_ sky130_fd_sc_hd__a22o_2
XFILLER_0_109_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17894_ VGND VPWR _03860_ _03794_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_205_500 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19633_ VGND VPWR VPWR VGND _05216_ _05052_ keymem.key_mem\[12\]\[109\] _05220_ sky130_fd_sc_hd__mux2_2
X_16845_ VGND VPWR _02986_ _09863_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_232_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_192_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_189_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16776_ VGND VPWR VGND VPWR _02923_ _02918_ _02917_ keylen _02922_ sky130_fd_sc_hd__o211ai_2
X_19564_ VGND VPWR VPWR VGND _05183_ _04992_ keymem.key_mem\[12\]\[76\] _05184_ sky130_fd_sc_hd__mux2_2
X_13988_ VPWR VGND VGND VPWR _09383_ _09460_ _09349_ sky130_fd_sc_hd__nor2_2
X_15727_ enc_block.sword_ctr_reg\[1\] _11183_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[23\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_18515_ VPWR VGND VPWR VGND _04395_ _04318_ _04393_ sky130_fd_sc_hd__or2_2
XFILLER_0_232_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12939_ VPWR VGND VPWR VGND _08464_ keymem.key_mem\[6\]\[77\] _07760_ keymem.key_mem\[11\]\[77\]
+ _07838_ _08465_ sky130_fd_sc_hd__a221o_2
XFILLER_0_5_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19495_ VGND VPWR VPWR VGND _05138_ _04943_ keymem.key_mem\[12\]\[44\] _05147_ sky130_fd_sc_hd__mux2_2
XFILLER_0_34_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_87_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_29_811 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15658_ VPWR VGND VPWR VGND _11114_ _11063_ _11115_ _10872_ _10997_ sky130_fd_sc_hd__or4b_2
XFILLER_0_47_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18446_ VGND VPWR _04332_ enc_block.block_w1_reg\[26\] enc_block.block_w0_reg\[1\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_238_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14609_ VGND VPWR VGND VPWR _10076_ _10032_ keymem.prev_key0_reg\[100\] _10077_ sky130_fd_sc_hd__a21o_2
X_18377_ VGND VPWR VGND VPWR _04270_ _04269_ _04271_ _03966_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_111_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_200_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15589_ VPWR VGND VPWR VGND _11047_ _11045_ _11046_ sky130_fd_sc_hd__or2_2
XFILLER_0_145_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_51_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17328_ VGND VPWR VGND VPWR _02750_ keymem.prev_key0_reg\[91\] _02864_ _03421_ sky130_fd_sc_hd__a21o_2
XFILLER_0_70_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17259_ _02460_ _03359_ keymem.prev_key0_reg\[84\] _02461_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_20270_ VGND VPWR VPWR VGND _05558_ _02608_ keymem.key_mem\[9\]\[22\] _05560_ sky130_fd_sc_hd__mux2_2
XFILLER_0_59_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_1017 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_216_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23960_ VGND VPWR VPWR VGND clk _00453_ reset_n keymem.key_mem\[13\]\[81\] sky130_fd_sc_hd__dfrtp_2
X_22911_ VGND VPWR VGND VPWR _06912_ _11559_ _03860_ _06884_ _02338_ sky130_fd_sc_hd__a211o_2
XFILLER_0_166_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23891_ VGND VPWR VPWR VGND clk _00384_ reset_n keymem.key_mem\[13\]\[12\] sky130_fd_sc_hd__dfrtp_2
X_25630_ VGND VPWR VPWR VGND clk _02123_ reset_n keymem.key_mem\[0\]\[87\] sky130_fd_sc_hd__dfrtp_2
X_22842_ VPWR VGND VPWR VGND _06870_ keymem.rcon_reg\[3\] keymem.rcon_logic.tmp_rcon\[0\]
+ sky130_fd_sc_hd__or2_2
XFILLER_0_195_215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_78_243 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25561_ VGND VPWR VPWR VGND clk _02054_ reset_n keymem.key_mem\[0\]\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22773_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[84\] _06837_ _06836_ _05006_ _02120_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_195_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_52_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24512_ VGND VPWR VPWR VGND clk _01005_ reset_n keymem.key_mem\[9\]\[121\] sky130_fd_sc_hd__dfrtp_2
X_21724_ VGND VPWR VPWR VGND _06330_ _03193_ keymem.key_mem\[4\]\[64\] _06332_ sky130_fd_sc_hd__mux2_2
XFILLER_0_52_1157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25492_ VGND VPWR VPWR VGND clk _01985_ reset_n keymem.key_mem\[1\]\[77\] sky130_fd_sc_hd__dfrtp_2
X_24443_ VGND VPWR VPWR VGND clk _00936_ reset_n keymem.key_mem\[9\]\[52\] sky130_fd_sc_hd__dfrtp_2
X_21655_ VGND VPWR _01555_ _06295_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20606_ VGND VPWR VPWR VGND _05736_ _03082_ keymem.key_mem\[8\]\[53\] _05737_ sky130_fd_sc_hd__mux2_2
XFILLER_0_266_1158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24374_ VGND VPWR VPWR VGND clk _00867_ reset_n keymem.key_mem\[10\]\[111\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_30_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21586_ VGND VPWR _06258_ _06257_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_793 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23325_ VPWR VGND _07204_ enc_block.block_w1_reg\[15\] enc_block.block_w1_reg\[11\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_20537_ VGND VPWR _01032_ _05700_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_144_392 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23256_ VGND VPWR _07142_ enc_block.block_w2_reg\[4\] _07141_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20468_ VGND VPWR _01000_ _05663_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_162_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22207_ VGND VPWR VPWR VGND _06589_ _02873_ keymem.key_mem\[2\]\[32\] _06591_ sky130_fd_sc_hd__mux2_2
XFILLER_0_242_1180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20399_ VGND VPWR _05627_ _05533_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23187_ VGND VPWR VPWR VGND _06880_ _07080_ keymem.prev_key1_reg\[125\] _07081_ sky130_fd_sc_hd__mux2_2
XFILLER_0_219_625 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_203_1142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22138_ VGND VPWR _06554_ _06553_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_218_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_246_455 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14960_ VGND VPWR VGND VPWR _10424_ _10423_ _10422_ keymem.prev_key1_reg\[13\] _09003_
+ _09002_ sky130_fd_sc_hd__a32o_2
X_22069_ VGND VPWR VPWR VGND _06516_ _05024_ keymem.key_mem\[3\]\[96\] _06517_ sky130_fd_sc_hd__mux2_2
X_13911_ VGND VPWR _09383_ _09382_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_227_691 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14891_ VPWR VGND VGND VPWR _10223_ _09690_ _10354_ _10355_ _10356_ sky130_fd_sc_hd__and4b_2
XFILLER_0_261_458 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16630_ VPWR VGND VPWR VGND _02785_ _02677_ _02775_ key[156] _02723_ _02786_ sky130_fd_sc_hd__a221o_2
X_13842_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[25\] _08956_ _09314_ _08943_ _09264_
+ _09265_ sky130_fd_sc_hd__a32oi_2
X_25828_ VGND VPWR VPWR VGND clk _02321_ reset_n enc_block.block_w3_reg\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_69_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_226_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_251_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_202_536 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16561_ VGND VPWR VGND VPWR _02720_ _11151_ key[153] _02707_ _02719_ sky130_fd_sc_hd__a211o_2
X_13773_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[24\] _08956_ _09245_ _08943_ _09243_
+ _09244_ sky130_fd_sc_hd__a32oi_2
X_25759_ keymem.prev_key1_reg\[75\] clk _02252_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_18300_ VPWR VGND VGND VPWR _04201_ _04202_ _04190_ sky130_fd_sc_hd__nor2_2
X_15512_ VGND VPWR VGND VPWR _10972_ _10971_ _10970_ _09868_ sky130_fd_sc_hd__o21a_2
X_19280_ VPWR VGND keymem.key_mem_we _05015_ _03409_ VPWR VGND sky130_fd_sc_hd__and2_2
X_12724_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[56\] _07843_ keymem.key_mem\[12\]\[56\]
+ _07620_ _08271_ sky130_fd_sc_hd__a22o_2
X_16492_ VPWR VGND VPWR VGND _02653_ keymem.prev_key1_reg\[87\] sky130_fd_sc_hd__inv_2
XFILLER_0_139_142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_151_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18231_ VGND VPWR _04138_ _03947_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_242_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15443_ VGND VPWR VGND VPWR _09981_ keymem.prev_key1_reg\[107\] _10904_ _09941_ sky130_fd_sc_hd__nand3_2
X_12655_ VGND VPWR VGND VPWR _08209_ _08008_ keymem.key_mem\[2\]\[49\] _08206_ _08208_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_84_279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18162_ VGND VPWR VGND VPWR _04072_ _03951_ _04075_ _00282_ sky130_fd_sc_hd__a21o_2
X_15374_ VGND VPWR _10836_ _10835_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12586_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[43\] _07845_ keymem.key_mem\[1\]\[43\]
+ _07901_ _08146_ sky130_fd_sc_hd__a22o_2
XFILLER_0_26_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_655 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17113_ VGND VPWR _03228_ _09541_ _00080_ _03227_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_14325_ VGND VPWR _09795_ _08935_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_25_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18093_ VPWR VGND _04012_ enc_block.block_w3_reg\[7\] enc_block.block_w3_reg\[2\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_52_165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_1397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17044_ VGND VPWR VPWR VGND _03164_ _03165_ _11624_ _03166_ sky130_fd_sc_hd__or3_2
X_14256_ VGND VPWR _00013_ _09726_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13207_ VGND VPWR VGND VPWR _08706_ _07968_ keymem.key_mem\[9\]\[104\] _08705_ _07574_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_110_226 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14187_ VGND VPWR _09658_ _09217_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_110_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13138_ VPWR VGND VPWR VGND _08643_ keymem.key_mem\[11\]\[97\] _07781_ keymem.key_mem\[10\]\[97\]
+ _07865_ _08644_ sky130_fd_sc_hd__a221o_2
X_18995_ _04824_ _04826_ _04560_ _04825_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_252_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13069_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[90\] _07722_ keymem.key_mem\[2\]\[90\]
+ _08131_ _08582_ sky130_fd_sc_hd__a22o_2
XFILLER_0_188_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17946_ VGND VPWR VGND VPWR _03670_ keymem.prev_key1_reg\[106\] _03530_ _03895_ sky130_fd_sc_hd__a21o_2
X_17877_ VGND VPWR VGND VPWR _03670_ keymem.prev_key1_reg\[84\] _03362_ _03848_ sky130_fd_sc_hd__a21o_2
XFILLER_0_206_864 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19616_ VGND VPWR VPWR VGND _05205_ _05035_ keymem.key_mem\[12\]\[101\] _05211_ sky130_fd_sc_hd__mux2_2
X_16828_ VGND VPWR VGND VPWR _10828_ _11456_ _02970_ _02969_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_75_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_221_834 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_49_906 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19547_ VPWR VGND VGND VPWR _05175_ keymem.key_mem\[12\]\[68\] _05095_ sky130_fd_sc_hd__nand2_2
X_16759_ VGND VPWR VPWR VGND _02906_ _02907_ _10327_ _10080_ _10081_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_18_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_221_889 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19478_ VGND VPWR _05138_ _05091_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_64_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_580 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_152_54 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_267_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18429_ VGND VPWR _04316_ _04314_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_185_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_847 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_44_622 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21440_ VGND VPWR _01454_ _06181_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_90_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_228_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_12_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_666 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21371_ VGND VPWR _01421_ _06145_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_160_126 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_86_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20322_ VGND VPWR VPWR VGND _05580_ _03025_ keymem.key_mem\[9\]\[47\] _05587_ sky130_fd_sc_hd__mux2_2
X_23110_ VGND VPWR _02272_ _07033_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_128_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_198 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24090_ VGND VPWR VPWR VGND clk _00583_ reset_n keymem.key_mem\[12\]\[83\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_40_850 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20253_ VGND VPWR VPWR VGND _05546_ _11099_ keymem.key_mem\[9\]\[14\] _05551_ sky130_fd_sc_hd__mux2_2
X_23041_ VGND VPWR _02245_ _06991_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_12_574 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20184_ VGND VPWR _00867_ _05512_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_239_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24992_ VGND VPWR VPWR VGND clk _01485_ reset_n keymem.key_mem\[5\]\[89\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_23_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23943_ VGND VPWR VPWR VGND clk _00436_ reset_n keymem.key_mem\[13\]\[64\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_239_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_93_1246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_252_981 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23874_ VGND VPWR VPWR VGND clk _00367_ reset_n enc_block.block_w2_reg\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_174_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_93_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25613_ VGND VPWR VPWR VGND clk _02106_ reset_n keymem.key_mem\[0\]\[70\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_223_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22825_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[124\] _06839_ _03864_ _05083_ _02160_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_6_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1168 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_196_579 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25544_ VGND VPWR VPWR VGND clk _02037_ reset_n keymem.key_mem\[0\]\[1\] sky130_fd_sc_hd__dfrtp_2
X_22756_ VGND VPWR VPWR VGND _06833_ keymem.key_mem\[0\]\[73\] _03268_ _06843_ sky130_fd_sc_hd__mux2_2
XFILLER_0_211_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21707_ VGND VPWR VPWR VGND _06319_ _03108_ keymem.key_mem\[4\]\[56\] _06323_ sky130_fd_sc_hd__mux2_2
XFILLER_0_109_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25475_ VGND VPWR VPWR VGND clk _01968_ reset_n keymem.key_mem\[1\]\[60\] sky130_fd_sc_hd__dfrtp_2
X_22687_ VGND VPWR _02067_ _06815_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_30_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24426_ VGND VPWR VPWR VGND clk _00919_ reset_n keymem.key_mem\[9\]\[35\] sky130_fd_sc_hd__dfrtp_2
X_12440_ VGND VPWR VGND VPWR _08014_ _08008_ keymem.key_mem\[2\]\[29\] _08010_ _08013_
+ sky130_fd_sc_hd__a211o_2
X_21638_ VGND VPWR VPWR VGND _06286_ _02660_ keymem.key_mem\[4\]\[23\] _06287_ sky130_fd_sc_hd__mux2_2
XFILLER_0_63_953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_370 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_168_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24357_ VGND VPWR VPWR VGND clk _00850_ reset_n keymem.key_mem\[10\]\[94\] sky130_fd_sc_hd__dfrtp_2
X_12371_ VGND VPWR VGND VPWR _07547_ keymem.key_mem\[2\]\[23\] _07947_ _07949_ _07951_
+ _07950_ sky130_fd_sc_hd__a2111o_2
X_21569_ VGND VPWR VPWR VGND _06242_ _03620_ keymem.key_mem\[5\]\[120\] _06249_ sky130_fd_sc_hd__mux2_2
XFILLER_0_151_137 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_34_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14110_ VGND VPWR VGND VPWR _09407_ _09479_ _09581_ _09380_ sky130_fd_sc_hd__a21oi_2
X_23308_ VPWR VGND VPWR VGND block[10] _03979_ enc_block.block_w1_reg\[10\] _03977_
+ _07189_ sky130_fd_sc_hd__a22o_2
X_15090_ VGND VPWR VGND VPWR _10554_ _10500_ _10472_ _10463_ _10464_ sky130_fd_sc_hd__a211o_2
XFILLER_0_65_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24288_ VGND VPWR VPWR VGND clk _00781_ reset_n keymem.key_mem\[10\]\[25\] sky130_fd_sc_hd__dfrtp_2
X_14041_ VGND VPWR _09513_ _09512_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_31_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23239_ VPWR VGND VGND VPWR _07126_ _07127_ _04019_ sky130_fd_sc_hd__nor2_2
XFILLER_0_24_1012 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17800_ VPWR VGND VPWR VGND _03127_ _03796_ keymem.prev_key0_reg\[58\] _03788_ _00199_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_101_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_712 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_219_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18780_ VPWR VGND _04633_ _04632_ enc_block.round_key\[35\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_247_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15992_ VGND VPWR VPWR VGND _11041_ keymem.key_mem\[14\]\[16\] _11447_ _11448_ sky130_fd_sc_hd__mux2_2
XFILLER_0_98_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14943_ VPWR VGND VPWR VGND _10407_ enc_block.block_w0_reg\[11\] _09273_ sky130_fd_sc_hd__or2_2
XFILLER_0_101_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17731_ VGND VPWR _00173_ _03753_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_190_1_Right_791 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_175_1336 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14874_ VPWR VGND VPWR VGND _10196_ _10338_ _10339_ _09207_ _09944_ sky130_fd_sc_hd__or4b_2
X_17662_ VGND VPWR _00153_ _03704_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_251_1213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_202_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_72_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1344 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19401_ VGND VPWR VGND VPWR _05096_ keymem.key_mem_we _09537_ _05093_ _00500_ sky130_fd_sc_hd__a31o_2
X_13825_ VGND VPWR _09297_ _09296_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16613_ VGND VPWR VGND VPWR _10075_ _10056_ _02769_ _09240_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_76_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17593_ VPWR VGND VGND VPWR _11456_ _03652_ key[253] sky130_fd_sc_hd__nor2_2
X_19332_ VGND VPWR VPWR VGND _05046_ _05048_ keymem.key_mem\[13\]\[107\] _05049_ sky130_fd_sc_hd__mux2_2
X_16544_ VGND VPWR _02703_ keymem.prev_key0_reg\[57\] keymem.prev_key0_reg\[89\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
X_13756_ VPWR VGND VGND VPWR _09228_ _09051_ _09086_ sky130_fd_sc_hd__nand2_2
XFILLER_0_97_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_31_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_57_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12707_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[54\] _08216_ keymem.key_mem\[6\]\[54\]
+ _07711_ _08256_ sky130_fd_sc_hd__a22o_2
X_16475_ VPWR VGND VPWR VGND _02631_ _02635_ _02636_ _02625_ _02630_ sky130_fd_sc_hd__or4b_2
X_19263_ VGND VPWR VGND VPWR _05004_ keymem.key_mem_we _03347_ _04999_ _00454_ sky130_fd_sc_hd__a31o_2
XFILLER_0_167_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13687_ VPWR VGND VPWR VGND _09031_ _09065_ _08971_ _08957_ _09159_ sky130_fd_sc_hd__or4_2
XFILLER_0_186_1410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15426_ VGND VPWR VGND VPWR _10519_ _10682_ _10887_ _10575_ sky130_fd_sc_hd__a21oi_2
X_18214_ VPWR VGND VPWR VGND _04122_ block[109] _03959_ enc_block.block_w2_reg\[13\]
+ _03954_ _04123_ sky130_fd_sc_hd__a221o_2
XFILLER_0_112_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19194_ VPWR VGND keymem.key_mem_we _04963_ _03099_ VPWR VGND sky130_fd_sc_hd__and2_2
X_12638_ VGND VPWR _08193_ _07560_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_108_1_Left_375 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_527 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_666 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18145_ VPWR VGND VPWR VGND _04059_ block[103] _03980_ enc_block.block_w3_reg\[7\]
+ _04007_ _04060_ sky130_fd_sc_hd__a221o_2
XFILLER_0_186_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15357_ VPWR VGND _10819_ keymem.prev_key0_reg\[74\] keymem.prev_key0_reg\[42\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
X_12569_ VGND VPWR _08131_ _07732_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14308_ VPWR VGND VPWR VGND _09591_ _09777_ _09617_ _09776_ _09778_ sky130_fd_sc_hd__or4_2
XFILLER_0_103_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18076_ VGND VPWR _03996_ enc_block.block_w2_reg\[10\] enc_block.block_w1_reg\[18\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_700 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15288_ VPWR VGND VPWR VGND _10749_ _10541_ _10498_ _10528_ _10750_ sky130_fd_sc_hd__a22o_2
XFILLER_0_41_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_40_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_83_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17027_ VGND VPWR VPWR VGND _03084_ keymem.key_mem\[14\]\[60\] _03150_ _03151_ sky130_fd_sc_hd__mux2_2
X_14239_ VGND VPWR VGND VPWR _09709_ _09639_ _09710_ keymem.prev_key0_reg\[97\] sky130_fd_sc_hd__a21oi_2
XFILLER_0_262_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_894 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_123_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_7_Right_7 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18978_ VPWR VGND VGND VPWR _04810_ _04811_ _04382_ sky130_fd_sc_hd__nor2_2
XFILLER_0_197_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17929_ VGND VPWR VPWR VGND _03874_ _03883_ keymem.prev_key0_reg\[100\] _03884_ sky130_fd_sc_hd__mux2_2
XFILLER_0_20_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_193_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20940_ VPWR VGND keymem.key_mem\[7\]\[79\] _05917_ _05899_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_234_1411 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20871_ VGND VPWR VGND VPWR _05879_ keymem.key_mem_we _03025_ _05864_ _01187_ sky130_fd_sc_hd__a31o_2
XFILLER_0_191_1182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_234_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22610_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[120\] _06777_ _06776_ _05075_ _02028_
+ sky130_fd_sc_hd__a22o_2
X_23590_ VGND VPWR VPWR VGND clk _00091_ reset_n keymem.key_mem\[14\]\[79\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_822 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_130_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22541_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[70\] _06754_ _06753_ _04983_ _01978_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_9_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25260_ VGND VPWR VPWR VGND clk _01753_ reset_n keymem.key_mem\[3\]\[101\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_8_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22472_ VGND VPWR _01937_ _06730_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_45_953 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_63_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24211_ VGND VPWR VPWR VGND clk _00704_ reset_n keymem.key_mem\[11\]\[76\] sky130_fd_sc_hd__dfrtp_2
X_21423_ VGND VPWR _01446_ _06172_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_165_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25191_ VGND VPWR VPWR VGND clk _01684_ reset_n keymem.key_mem\[3\]\[32\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_31_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24142_ VGND VPWR VPWR VGND clk _00635_ reset_n keymem.key_mem\[11\]\[7\] sky130_fd_sc_hd__dfrtp_2
X_21354_ VGND VPWR _01413_ _06136_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_32_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20305_ VGND VPWR VPWR VGND _05569_ _02945_ keymem.key_mem\[9\]\[39\] _05578_ sky130_fd_sc_hd__mux2_2
X_24073_ VGND VPWR VPWR VGND clk _00566_ reset_n keymem.key_mem\[12\]\[66\] sky130_fd_sc_hd__dfrtp_2
X_21285_ VGND VPWR VPWR VGND _06098_ _03580_ keymem.key_mem\[6\]\[114\] _06099_ sky130_fd_sc_hd__mux2_2
XFILLER_0_97_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23024_ VGND VPWR VPWR VGND _02238_ _03155_ _03160_ _06925_ _06981_ sky130_fd_sc_hd__o31a_2
X_20236_ VGND VPWR VPWR VGND _05535_ _10284_ keymem.key_mem\[9\]\[6\] _05542_ sky130_fd_sc_hd__mux2_2
XFILLER_0_204_1270 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20167_ VGND VPWR _00859_ _05503_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_102_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_122_2_Left_593 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_217_948 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_200_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20098_ VGND VPWR _00826_ _05467_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24975_ VGND VPWR VPWR VGND clk _01468_ reset_n keymem.key_mem\[5\]\[72\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23926_ VGND VPWR VPWR VGND clk _00419_ reset_n keymem.key_mem\[13\]\[47\] sky130_fd_sc_hd__dfrtp_2
X_11940_ VGND VPWR VGND VPWR _07525_ _07543_ _07526_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_252_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_196_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11871_ VGND VPWR result[102] _07499_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23857_ VGND VPWR VPWR VGND clk _00350_ reset_n enc_block.block_w2_reg\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_170_1222 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_19_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_1049 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_252_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13610_ VGND VPWR _09082_ _09081_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_79_371 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22808_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[109\] _06858_ _06857_ _05052_ _02145_
+ sky130_fd_sc_hd__a22o_2
X_14590_ VGND VPWR VGND VPWR _09559_ _09386_ _09480_ _09419_ _10058_ sky130_fd_sc_hd__o22a_2
XFILLER_0_79_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23788_ VGND VPWR VPWR VGND clk _00281_ reset_n enc_block.block_w0_reg\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13541_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[6\] _08989_ _09013_ _08983_ _08980_
+ _08981_ sky130_fd_sc_hd__a32oi_2
X_25527_ VGND VPWR VPWR VGND clk _02020_ reset_n keymem.key_mem\[1\]\[112\] sky130_fd_sc_hd__dfrtp_2
X_22739_ VGND VPWR VPWR VGND _06833_ keymem.key_mem\[0\]\[64\] _03194_ _06835_ sky130_fd_sc_hd__mux2_2
XFILLER_0_149_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16260_ VPWR VGND VGND VPWR _11473_ _02424_ _11182_ sky130_fd_sc_hd__nor2_2
X_13472_ VPWR VGND VPWR VGND _08944_ enc_block.sword_ctr_reg\[0\] sky130_fd_sc_hd__inv_2
X_25458_ VGND VPWR VPWR VGND clk _01951_ reset_n keymem.key_mem\[1\]\[43\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_109_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15211_ VPWR VGND VGND VPWR _10535_ _10674_ _10633_ sky130_fd_sc_hd__nor2_2
XFILLER_0_36_975 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12423_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[28\] _07587_ keymem.key_mem\[11\]\[28\]
+ _07600_ _07998_ sky130_fd_sc_hd__a22o_2
X_24409_ VGND VPWR VPWR VGND clk _00902_ reset_n keymem.key_mem\[9\]\[18\] sky130_fd_sc_hd__dfrtp_2
X_16191_ VGND VPWR VGND VPWR _02356_ _11348_ _11292_ _11371_ _11506_ sky130_fd_sc_hd__a211o_2
X_25389_ VGND VPWR VPWR VGND clk _01882_ reset_n keymem.key_mem\[2\]\[102\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_129_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15142_ VPWR VGND VPWR VGND _10599_ _10605_ _10600_ _10598_ _10606_ sky130_fd_sc_hd__or4_2
X_12354_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[22\] _07596_ keymem.key_mem\[8\]\[22\]
+ _07752_ _07935_ sky130_fd_sc_hd__a22o_2
XFILLER_0_65_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_105_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15073_ VPWR VGND VGND VPWR _10536_ _10537_ _10489_ sky130_fd_sc_hd__nor2_2
XFILLER_0_50_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_120_321 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_266_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19950_ VGND VPWR VPWR VGND _05389_ _09537_ keymem.key_mem\[10\]\[0\] _05390_ sky130_fd_sc_hd__mux2_2
XFILLER_0_120_332 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12285_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[17\] _07695_ keymem.key_mem\[14\]\[17\]
+ _07782_ _07871_ sky130_fd_sc_hd__a22o_2
X_14024_ VGND VPWR VGND VPWR _09494_ _09389_ _09496_ _09495_ sky130_fd_sc_hd__a21oi_2
X_18901_ VPWR VGND _04742_ _04741_ enc_block.round_key\[47\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_19881_ VGND VPWR VPWR VGND _05350_ keymem.key_mem\[11\]\[97\] _03474_ _05352_ sky130_fd_sc_hd__mux2_2
XFILLER_0_120_387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_248_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18832_ VPWR VGND VPWR VGND _04680_ enc_block.round_key\[40\] _04679_ sky130_fd_sc_hd__or2_2
X_18763_ VGND VPWR _04617_ enc_block.block_w1_reg\[1\] _04616_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15975_ VPWR VGND VPWR VGND _11428_ _11430_ _11429_ _11425_ _11431_ sky130_fd_sc_hd__or4_2
XFILLER_0_223_918 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_191_1_Right_792 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17714_ VPWR VGND VPWR VGND _02740_ _03742_ keymem.prev_key0_reg\[26\] _03730_ _00167_
+ sky130_fd_sc_hd__a22o_2
X_14926_ VGND VPWR VGND VPWR enc_block.block_w2_reg\[9\] _09269_ _10387_ _10388_ _10390_
+ _10389_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_262_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1166 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18694_ VPWR VGND VPWR VGND _04555_ _04341_ _04553_ sky130_fd_sc_hd__or2_2
XFILLER_0_117_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_251_1032 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17645_ VGND VPWR VPWR VGND _03681_ _03692_ keymem.prev_key0_reg\[7\] _03693_ sky130_fd_sc_hd__mux2_2
X_14857_ VGND VPWR _10322_ _09729_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_202_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_37_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_472 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13808_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[30\] _08969_ _09280_ _08964_ _09278_
+ _09279_ sky130_fd_sc_hd__a32oi_2
X_14788_ VGND VPWR VGND VPWR _09348_ _09352_ _09335_ _09486_ _10254_ sky130_fd_sc_hd__o22a_2
X_17576_ VPWR VGND VGND VPWR _03637_ _02755_ _02756_ sky130_fd_sc_hd__nand2_2
X_19315_ VPWR VGND keymem.key_mem_we _05037_ _03506_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13739_ VGND VPWR _09211_ _09210_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16527_ VPWR VGND VPWR VGND _02687_ _10086_ _02684_ _02685_ _02686_ _10096_ sky130_fd_sc_hd__o311a_2
XFILLER_0_42_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_599 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_220_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19246_ VGND VPWR VPWR VGND _04993_ _04992_ keymem.key_mem\[13\]\[76\] _04994_ sky130_fd_sc_hd__mux2_2
XFILLER_0_229_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16458_ VPWR VGND VPWR VGND _02618_ _11477_ _11486_ _11323_ _02378_ _02619_ sky130_fd_sc_hd__a221o_2
XFILLER_0_45_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15409_ VGND VPWR VGND VPWR _10528_ _10538_ _10870_ _10546_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_6_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19177_ VGND VPWR _00420_ _04952_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16389_ VGND VPWR _00033_ _02551_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_147_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18128_ VPWR VGND _04044_ enc_block.block_w1_reg\[22\] enc_block.block_w2_reg\[14\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_83_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_147_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_444 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_48_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_83_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18059_ VGND VPWR _03980_ _03979_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21070_ VGND VPWR _05986_ _10913_ _01279_ _05985_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_1_585 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20021_ VGND VPWR _00789_ _05427_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_158_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24760_ VGND VPWR VPWR VGND clk _01253_ reset_n keymem.key_mem\[7\]\[113\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_158_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21972_ VGND VPWR _01702_ _06465_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_94_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_154_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23711_ keymem.prev_key0_reg\[67\] clk _00208_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_174_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20923_ VGND VPWR VGND VPWR _05907_ keymem.key_mem_we _03252_ _05893_ _01211_ sky130_fd_sc_hd__a31o_2
XFILLER_0_7_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24691_ VGND VPWR VPWR VGND clk _01184_ reset_n keymem.key_mem\[7\]\[44\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23642_ VGND VPWR VPWR VGND clk _00002_ reset_n keymem.round_ctr_rst sky130_fd_sc_hd__dfrtp_2
XFILLER_0_7_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20854_ VGND VPWR VPWR VGND _05867_ _04933_ keymem.key_mem\[7\]\[39\] _05871_ sky130_fd_sc_hd__mux2_2
XFILLER_0_193_302 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_238_Right_107 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_717 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_7_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23573_ VGND VPWR VPWR VGND clk _00074_ reset_n keymem.key_mem\[14\]\[62\] sky130_fd_sc_hd__dfrtp_2
X_20785_ VGND VPWR _01147_ _05833_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25312_ VGND VPWR VPWR VGND clk _01805_ reset_n keymem.key_mem\[2\]\[25\] sky130_fd_sc_hd__dfrtp_2
X_22524_ VGND VPWR _01970_ _06749_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_9_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25243_ VGND VPWR VPWR VGND clk _01736_ reset_n keymem.key_mem\[3\]\[84\] sky130_fd_sc_hd__dfrtp_2
X_22455_ VGND VPWR _01929_ _06721_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_165_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1067 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21406_ VGND VPWR VPWR VGND _06162_ _02972_ keymem.key_mem\[5\]\[42\] _06164_ sky130_fd_sc_hd__mux2_2
XFILLER_0_66_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_126_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25174_ VGND VPWR VPWR VGND clk _01667_ reset_n keymem.key_mem\[3\]\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22386_ VGND VPWR _01897_ _06684_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_165_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24125_ VGND VPWR VPWR VGND clk _00618_ reset_n keymem.key_mem\[12\]\[118\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_66_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21337_ VGND VPWR _01405_ _06127_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_27_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_848 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_102_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24056_ VGND VPWR VPWR VGND clk _00549_ reset_n keymem.key_mem\[12\]\[49\] sky130_fd_sc_hd__dfrtp_2
X_12070_ VGND VPWR _07670_ _07556_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21268_ VGND VPWR VPWR VGND _06087_ _03533_ keymem.key_mem\[6\]\[106\] _06090_ sky130_fd_sc_hd__mux2_2
XFILLER_0_241_1289 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_229_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23007_ VGND VPWR _02231_ _06971_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20219_ VPWR VGND VPWR VGND _05240_ _05531_ _05530_ keymem.round_ctr_reg\[1\] sky130_fd_sc_hd__or3b_2
X_21199_ VGND VPWR VPWR VGND _06052_ _03267_ keymem.key_mem\[6\]\[73\] _06054_ sky130_fd_sc_hd__mux2_2
XFILLER_0_102_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15760_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[16\] _10402_ _11216_ _09255_ _11214_
+ _11215_ sky130_fd_sc_hd__a32oi_2
X_24958_ VGND VPWR VPWR VGND clk _01451_ reset_n keymem.key_mem\[5\]\[55\] sky130_fd_sc_hd__dfrtp_2
X_12972_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[80\] _07644_ _08494_ _08490_ _08495_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_176_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_172_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14711_ VPWR VGND VPWR VGND _10177_ _10178_ _10176_ _09798_ sky130_fd_sc_hd__or3b_2
X_11923_ VGND VPWR VPWR VGND encdec enc_block.round\[1\] dec_round_nr\[1\] _07526_
+ sky130_fd_sc_hd__mux2_2
X_15691_ VPWR VGND VPWR VGND _11147_ _09638_ _11108_ key[143] _11043_ _11148_ sky130_fd_sc_hd__a221o_2
X_23909_ VGND VPWR VPWR VGND clk _00402_ reset_n keymem.key_mem\[13\]\[30\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_73_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1352 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24889_ VGND VPWR VPWR VGND clk _01382_ reset_n keymem.key_mem\[6\]\[114\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_34_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14642_ VPWR VGND VGND VPWR _09362_ _09348_ _09440_ _10109_ sky130_fd_sc_hd__nor3_2
X_17430_ VGND VPWR VGND VPWR _03511_ _10838_ key[231] _03509_ _03510_ sky130_fd_sc_hd__a211o_2
X_11854_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[30\] dec_new_block\[94\]
+ _07491_ sky130_fd_sc_hd__mux2_2
XFILLER_0_200_623 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_197_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_77 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_196_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14573_ VPWR VGND VGND VPWR _10041_ _09907_ _09906_ sky130_fd_sc_hd__nand2_2
X_17361_ VGND VPWR VGND VPWR keylen _03451_ _03450_ _10323_ _02831_ _02832_ sky130_fd_sc_hd__a311oi_2
X_11785_ VGND VPWR result[59] _07456_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_94_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_103_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19100_ VPWR VGND keymem.key_mem\[13\]\[19\] _04905_ _04903_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_32_1166 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13524_ VPWR VGND VPWR VGND _08996_ enc_block.block_w0_reg\[4\] _08995_ sky130_fd_sc_hd__or2_2
X_16312_ VGND VPWR VPWR VGND _09927_ _02469_ key[148] _02476_ sky130_fd_sc_hd__mux2_2
X_17292_ VPWR VGND _03389_ _03388_ keymem.prev_key0_reg\[87\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_27_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_137_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_250_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19031_ VGND VPWR VGND VPWR _03958_ block[61] _04857_ _04858_ sky130_fd_sc_hd__a21o_2
X_16243_ VPWR VGND VGND VPWR _02406_ _02407_ _02405_ _02403_ _02408_ _09637_ sky130_fd_sc_hd__o221a_2
XFILLER_0_246_1123 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_187_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13455_ VGND VPWR _08927_ _08926_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_3_806 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_10_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12406_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[26\] _07644_ _07982_ _07978_ _07983_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_35_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16174_ VGND VPWR _02340_ _02339_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_10_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13386_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[122\] _07785_ keymem.key_mem\[2\]\[122\]
+ _08116_ _08867_ sky130_fd_sc_hd__a22o_2
XFILLER_0_144_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15125_ VGND VPWR VGND VPWR _10585_ _10583_ _10589_ _10588_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_80_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12337_ VPWR VGND VPWR VGND keymem.key_mem\[8\]\[20\] _07654_ keymem.key_mem\[1\]\[20\]
+ _07714_ _07920_ sky130_fd_sc_hd__a22o_2
XFILLER_0_45_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1192 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15056_ VGND VPWR _10520_ _10507_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_266_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19933_ VGND VPWR VPWR VGND _05372_ keymem.key_mem\[11\]\[122\] _03633_ _05379_ sky130_fd_sc_hd__mux2_2
X_12268_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[15\] _07724_ keymem.key_mem\[1\]\[15\]
+ _07855_ _07856_ sky130_fd_sc_hd__a22o_2
XFILLER_0_267_689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_208_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14007_ VGND VPWR VPWR VGND _09304_ _09246_ _09303_ _09479_ sky130_fd_sc_hd__or3_2
X_19864_ VGND VPWR VPWR VGND _05339_ keymem.key_mem\[11\]\[89\] _03409_ _05343_ sky130_fd_sc_hd__mux2_2
XFILLER_0_254_339 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12199_ VGND VPWR VGND VPWR _07792_ _07786_ keymem.key_mem\[10\]\[10\] _07789_ _07791_
+ sky130_fd_sc_hd__a211o_2
X_18815_ VPWR VGND VGND VPWR _04654_ _04665_ _04052_ sky130_fd_sc_hd__nor2_2
XFILLER_0_120_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19795_ VGND VPWR VPWR VGND _05303_ keymem.key_mem\[11\]\[56\] _03109_ _05307_ sky130_fd_sc_hd__mux2_2
XFILLER_0_170_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_207_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_155_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18746_ VGND VPWR VGND VPWR _04598_ _03951_ _04601_ _00340_ sky130_fd_sc_hd__a21o_2
XFILLER_0_194_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15958_ VPWR VGND VGND VPWR _11218_ _11257_ _11414_ _11308_ _11283_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_91_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_192_1_Right_793 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_155_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1022 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14909_ VGND VPWR VGND VPWR _09238_ _09165_ _10373_ keymem.prev_key1_reg\[104\] sky130_fd_sc_hd__a21oi_2
X_18677_ VPWR VGND VPWR VGND _04539_ block[89] _04487_ enc_block.block_w1_reg\[25\]
+ _04425_ _04540_ sky130_fd_sc_hd__a221o_2
XFILLER_0_235_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_210_409 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15889_ VGND VPWR _11345_ _11344_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_8_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17628_ VGND VPWR _03681_ _03674_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_8_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17559_ VPWR VGND VGND VPWR _03622_ _03240_ _02702_ sky130_fd_sc_hd__nand2_2
XFILLER_0_85_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_18_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20570_ VGND VPWR VPWR VGND _05714_ _02913_ keymem.key_mem\[8\]\[36\] _05718_ sky130_fd_sc_hd__mux2_2
XFILLER_0_229_1310 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_108_2_Right_180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19229_ VPWR VGND keymem.key_mem_we _04983_ _03245_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_5_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22240_ VGND VPWR VPWR VGND _06600_ _03035_ keymem.key_mem\[2\]\[48\] _06608_ sky130_fd_sc_hd__mux2_2
XFILLER_0_14_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_915 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_242_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_75_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22171_ VGND VPWR VPWR VGND _06565_ _11148_ keymem.key_mem\[2\]\[15\] _06572_ sky130_fd_sc_hd__mux2_2
XFILLER_0_203_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_242_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21122_ VGND VPWR _01304_ _06013_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_246_818 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_203_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_111_195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21053_ VGND VPWR VPWR VGND _05972_ _10098_ keymem.key_mem\[6\]\[4\] _05977_ sky130_fd_sc_hd__mux2_2
XFILLER_0_258_1049 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20004_ VGND VPWR _00781_ _05418_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_195_1339 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24812_ VGND VPWR VPWR VGND clk _01305_ reset_n keymem.key_mem\[6\]\[37\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_198_405 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25792_ keymem.prev_key1_reg\[108\] clk _02285_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_158_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1145 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24743_ VGND VPWR VPWR VGND clk _01236_ reset_n keymem.key_mem\[7\]\[96\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_94_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21955_ VGND VPWR _01694_ _06456_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_16_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20906_ VGND VPWR VGND VPWR _05898_ keymem.key_mem_we _03184_ _05893_ _01203_ sky130_fd_sc_hd__a31o_2
X_24674_ VGND VPWR VPWR VGND clk _01167_ reset_n keymem.key_mem\[7\]\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_222_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_1_Right_667 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21886_ VGND VPWR VPWR VGND _06403_ _04894_ keymem.key_mem\[3\]\[11\] _06419_ sky130_fd_sc_hd__mux2_2
XFILLER_0_210_954 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_210_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23625_ VGND VPWR VPWR VGND clk _00126_ reset_n keymem.key_mem\[14\]\[114\] sky130_fd_sc_hd__dfrtp_2
X_20837_ VGND VPWR VGND VPWR _05861_ keymem.key_mem_we _02862_ _05850_ _01171_ sky130_fd_sc_hd__a31o_2
XFILLER_0_49_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23556_ VGND VPWR VPWR VGND clk _00057_ reset_n keymem.key_mem\[14\]\[45\] sky130_fd_sc_hd__dfrtp_2
X_20768_ VGND VPWR _05824_ _05823_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22507_ VGND VPWR _01961_ _06741_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_181_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23487_ VPWR VGND VGND VPWR _07192_ _07349_ _04283_ sky130_fd_sc_hd__nor2_2
XFILLER_0_64_388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20699_ VGND VPWR _01109_ _05785_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_134_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25226_ VGND VPWR VPWR VGND clk _01719_ reset_n keymem.key_mem\[3\]\[67\] sky130_fd_sc_hd__dfrtp_2
X_13240_ VGND VPWR _08736_ _07746_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22438_ VGND VPWR _01921_ _06712_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_27_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13171_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[100\] _07799_ keymem.key_mem\[2\]\[100\]
+ _07546_ _08674_ sky130_fd_sc_hd__a22o_2
X_25157_ VGND VPWR VPWR VGND clk _01650_ reset_n keymem.key_mem\[4\]\[126\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22369_ VGND VPWR _01889_ _06675_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_66_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24108_ VGND VPWR VPWR VGND clk _00601_ reset_n keymem.key_mem\[12\]\[101\] sky130_fd_sc_hd__dfrtp_2
X_12122_ VPWR VGND VPWR VGND _07718_ keymem.key_mem\[9\]\[6\] _07717_ keymem.key_mem\[1\]\[6\]
+ _07715_ _07719_ sky130_fd_sc_hd__a221o_2
XFILLER_0_108_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_102_162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25088_ VGND VPWR VPWR VGND clk _01581_ reset_n keymem.key_mem\[4\]\[57\] sky130_fd_sc_hd__dfrtp_2
X_16930_ VGND VPWR VGND VPWR _02403_ _10278_ _03062_ _03063_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_248_188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24039_ VGND VPWR VPWR VGND clk _00532_ reset_n keymem.key_mem\[12\]\[32\] sky130_fd_sc_hd__dfrtp_2
X_12053_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[3\] _07652_ keymem.key_mem\[7\]\[3\]
+ _07650_ _07653_ sky130_fd_sc_hd__a22o_2
XFILLER_0_263_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_542 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16861_ VGND VPWR VGND VPWR _11025_ _11024_ _10386_ _03000_ sky130_fd_sc_hd__a21o_2
XFILLER_0_102_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18600_ VGND VPWR _04471_ enc_block.block_w3_reg\[9\] enc_block.block_w0_reg\[1\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15812_ VPWR VGND VGND VPWR _11267_ _11268_ _11262_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_117_1_Left_384 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19580_ VGND VPWR VGND VPWR _05192_ keymem.key_mem_we _03356_ _05187_ _00583_ sky130_fd_sc_hd__a31o_2
X_16792_ VGND VPWR VGND VPWR _02937_ _10732_ _10364_ _10363_ _10329_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_176_1272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_137_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1283 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18531_ VGND VPWR _04409_ enc_block.block_w0_reg\[2\] _04408_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15743_ VGND VPWR VGND VPWR _11199_ enc_block.block_w2_reg\[21\] enc_block.sword_ctr_reg\[1\]
+ enc_block.sword_ctr_reg\[0\] sky130_fd_sc_hd__and3b_2
XFILLER_0_99_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12955_ VPWR VGND VPWR VGND _08478_ keymem.key_mem\[1\]\[79\] _07715_ keymem.key_mem\[2\]\[79\]
+ _07698_ _08479_ sky130_fd_sc_hd__a221o_2
XFILLER_0_77_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_140 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11906_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[24\] dec_new_block\[120\]
+ _07517_ sky130_fd_sc_hd__mux2_2
XFILLER_0_73_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18462_ VPWR VGND VPWR VGND block[67] _03957_ enc_block.block_w0_reg\[3\] _03952_
+ _04347_ sky130_fd_sc_hd__a22o_2
XFILLER_0_90_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15674_ VGND VPWR VGND VPWR _10644_ _10528_ _10508_ _11131_ sky130_fd_sc_hd__a21o_2
X_12886_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[72\] _07579_ keymem.key_mem\[1\]\[72\]
+ _07800_ _08417_ sky130_fd_sc_hd__a22o_2
XFILLER_0_38_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_200_431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17413_ VPWR VGND VGND VPWR _03496_ key[229] _08929_ sky130_fd_sc_hd__nand2_2
X_11837_ VGND VPWR result[85] _07482_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14625_ VPWR VGND VGND VPWR _10093_ key[132] _10091_ sky130_fd_sc_hd__nand2_2
X_18393_ VGND VPWR _04285_ enc_block.block_w0_reg\[29\] _04214_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_536 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_157_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14556_ VPWR VGND VGND VPWR _09116_ _10024_ _09056_ sky130_fd_sc_hd__nor2_2
XFILLER_0_67_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17344_ VGND VPWR VPWR VGND _03384_ keymem.key_mem\[14\]\[92\] _03435_ _03436_ sky130_fd_sc_hd__mux2_2
X_11768_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[19\] dec_new_block\[51\]
+ _07448_ sky130_fd_sc_hd__mux2_2
X_13507_ enc_block.sword_ctr_reg\[1\] _08979_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[6\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_125_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14487_ VPWR VGND VPWR VGND _09955_ _09202_ _09680_ _09700_ _09956_ sky130_fd_sc_hd__or4bb_2
X_17275_ VPWR VGND VPWR VGND _03373_ _03370_ _03369_ key[213] _03366_ _03374_ sky130_fd_sc_hd__a221o_2
X_11699_ VGND VPWR result[16] _07413_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_10_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19014_ VPWR VGND VPWR VGND _04842_ block[59] _04837_ enc_block.block_w2_reg\[27\]
+ _04798_ _04843_ sky130_fd_sc_hd__a221o_2
XFILLER_0_109_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16226_ VPWR VGND VPWR VGND _02391_ _11338_ _11182_ _11205_ _02389_ _02390_ sky130_fd_sc_hd__o311a_2
X_13438_ VPWR VGND VPWR VGND _08913_ keymem.key_mem\[1\]\[127\] _07715_ keymem.key_mem\[2\]\[127\]
+ _07546_ _08914_ sky130_fd_sc_hd__a221o_2
XFILLER_0_148_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_915 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_45_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1276 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_144_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16157_ VPWR VGND VGND VPWR _11235_ _11611_ _11252_ sky130_fd_sc_hd__nor2_2
XFILLER_0_49_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13369_ VGND VPWR VGND VPWR _07780_ keymem.key_mem\[5\]\[120\] _08849_ _08851_ _08852_
+ _08736_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_12_959 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15108_ VGND VPWR _10572_ _10559_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16088_ VGND VPWR _11543_ _08935_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15039_ VPWR VGND VPWR VGND _10424_ _10445_ _10444_ _10419_ _10503_ sky130_fd_sc_hd__or4_2
X_19916_ VGND VPWR VPWR VGND _05361_ keymem.key_mem\[11\]\[114\] _03580_ _05370_ sky130_fd_sc_hd__mux2_2
XFILLER_0_20_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_840 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_259_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19847_ VGND VPWR VPWR VGND _05328_ keymem.key_mem\[11\]\[81\] _03339_ _05334_ sky130_fd_sc_hd__mux2_2
XFILLER_0_251_810 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1022 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19778_ VGND VPWR VPWR VGND _05292_ keymem.key_mem\[11\]\[48\] _03035_ _05298_ sky130_fd_sc_hd__mux2_2
XFILLER_0_64_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1139 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18729_ VPWR VGND VPWR VGND _04586_ _04443_ _04584_ sky130_fd_sc_hd__or2_2
XFILLER_0_91_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_578 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_155_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_193_1_Right_794 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21740_ VGND VPWR VPWR VGND _06330_ _03259_ keymem.key_mem\[4\]\[72\] _06340_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_175_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21671_ VGND VPWR VPWR VGND _06297_ _02945_ keymem.key_mem\[4\]\[39\] _06304_ sky130_fd_sc_hd__mux2_2
XFILLER_0_46_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_175_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23410_ VPWR VGND _07281_ _07280_ enc_block.round_key\[20\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_46_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_2_Left_550 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20622_ VGND VPWR VPWR VGND _05736_ _03161_ keymem.key_mem\[8\]\[61\] _05745_ sky130_fd_sc_hd__mux2_2
X_24390_ VGND VPWR VPWR VGND clk _00883_ reset_n keymem.key_mem\[10\]\[127\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_266_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_931 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_163_349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23341_ VPWR VGND _07219_ _07218_ enc_block.round_key\[13\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_116_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_34_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20553_ VGND VPWR VPWR VGND _05703_ _02786_ keymem.key_mem\[8\]\[28\] _05709_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_109_2_Right_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_127_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23272_ VPWR VGND VPWR VGND _07156_ _04874_ _07155_ enc_block.block_w3_reg\[6\] _07115_
+ _02311_ sky130_fd_sc_hd__a221o_2
XFILLER_0_85_1148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20484_ VGND VPWR _01008_ _05671_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_30_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25011_ VGND VPWR VPWR VGND clk _01504_ reset_n keymem.key_mem\[5\]\[108\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_171_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_28_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22223_ VGND VPWR VPWR VGND _06589_ _02955_ keymem.key_mem\[2\]\[40\] _06599_ sky130_fd_sc_hd__mux2_2
XFILLER_0_15_797 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_63_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_258_453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22154_ VGND VPWR _01787_ _06562_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_207_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21105_ VGND VPWR _01296_ _06004_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_182_1_Left_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22085_ VGND VPWR VPWR VGND _06516_ _05041_ keymem.key_mem\[3\]\[104\] _06525_ sky130_fd_sc_hd__mux2_2
X_21036_ VGND VPWR _01265_ _05966_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_103_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25775_ keymem.prev_key1_reg\[91\] clk _02268_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22987_ VGND VPWR _06960_ _06880_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12740_ VGND VPWR VGND VPWR _08286_ _07648_ keymem.key_mem\[2\]\[57\] _08285_ _07573_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_201_228 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_74_1575 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_96_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21938_ VGND VPWR VGND VPWR _06447_ keymem.key_mem_we _02894_ _06446_ _01686_ sky130_fd_sc_hd__a31o_2
X_24726_ VGND VPWR VPWR VGND clk _01219_ reset_n keymem.key_mem\[7\]\[79\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_215_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12671_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[51\] _07649_ keymem.key_mem\[4\]\[51\]
+ _07913_ _08223_ sky130_fd_sc_hd__a22o_2
X_24657_ VGND VPWR VPWR VGND clk _01150_ reset_n keymem.key_mem\[7\]\[10\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_67_1_Right_668 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_210_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21869_ VPWR VGND keymem.key_mem\[3\]\[3\] _06410_ _06406_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_249_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_214_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14410_ VPWR VGND VGND VPWR _09879_ _09487_ _09450_ sky130_fd_sc_hd__nand2_2
XFILLER_0_38_856 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23608_ VGND VPWR VPWR VGND clk _00109_ reset_n keymem.key_mem\[14\]\[97\] sky130_fd_sc_hd__dfrtp_2
X_15390_ VPWR VGND VGND VPWR _10511_ _10851_ _10627_ sky130_fd_sc_hd__nor2_2
X_24588_ VGND VPWR VPWR VGND clk _01081_ reset_n keymem.key_mem\[8\]\[69\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_64_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_249_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14341_ VGND VPWR VGND VPWR _09221_ _08999_ _09097_ _09157_ _09811_ sky130_fd_sc_hd__o22a_2
XFILLER_0_64_152 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_110_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23539_ VGND VPWR VPWR VGND clk _00040_ reset_n keymem.key_mem\[14\]\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_231_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17060_ VPWR VGND VPWR VGND _03181_ key[191] _10322_ sky130_fd_sc_hd__or2_2
XFILLER_0_11_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14272_ VPWR VGND VPWR VGND _09742_ _09480_ _09305_ sky130_fd_sc_hd__or2_2
XFILLER_0_145_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16011_ VGND VPWR _11466_ _11465_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_33_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25209_ VGND VPWR VPWR VGND clk _01702_ reset_n keymem.key_mem\[3\]\[50\] sky130_fd_sc_hd__dfrtp_2
X_13223_ VPWR VGND VPWR VGND _08720_ keymem.key_mem\[3\]\[105\] _08009_ keymem.key_mem\[14\]\[105\]
+ _07963_ _08721_ sky130_fd_sc_hd__a221o_2
XFILLER_0_145_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_572 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_723 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1054 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_265_902 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13154_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[98\] _08577_ _08658_ _08654_ _08659_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_20_244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_237_626 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12105_ VGND VPWR _07703_ _07702_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_221_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1210 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13085_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[92\] _07834_ keymem.key_mem\[11\]\[92\]
+ _07809_ _08596_ sky130_fd_sc_hd__a22o_2
X_17962_ VGND VPWR VPWR VGND _03876_ key[239] keymem.prev_key1_reg\[111\] _03906_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_40_1232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19701_ VGND VPWR _05257_ _10913_ _00639_ _05243_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_256_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16913_ VGND VPWR _00061_ _03047_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12036_ VGND VPWR _07637_ _07636_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_178_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_256_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17893_ VGND VPWR _03859_ _02947_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_254_1200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19632_ VGND VPWR _00608_ _05219_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16844_ VPWR VGND VPWR VGND _02984_ _10902_ _02977_ key[171] _02875_ _02985_ sky130_fd_sc_hd__a221o_2
XFILLER_0_217_383 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_256_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19563_ VGND VPWR _05183_ _05091_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_189_246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16775_ VGND VPWR VGND VPWR _02922_ _02919_ _10146_ _02920_ _02921_ sky130_fd_sc_hd__a211o_2
XFILLER_0_152_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13987_ VPWR VGND VGND VPWR _09396_ _09459_ _09349_ sky130_fd_sc_hd__nor2_2
XFILLER_0_205_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1288 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18514_ VPWR VGND VGND VPWR _04394_ _04318_ _04393_ sky130_fd_sc_hd__nand2_2
X_15726_ VGND VPWR _11182_ _11181_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_125_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19494_ VGND VPWR _00543_ _05146_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12938_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[77\] _07587_ keymem.key_mem\[12\]\[77\]
+ _07621_ _08464_ sky130_fd_sc_hd__a22o_2
XFILLER_0_232_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18445_ VPWR VGND _04331_ enc_block.block_w2_reg\[18\] enc_block.block_w3_reg\[10\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_87_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15657_ VPWR VGND VGND VPWR _10485_ _10646_ _10672_ _11114_ sky130_fd_sc_hd__nor3_2
XFILLER_0_28_300 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_29_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12869_ VPWR VGND VPWR VGND _08401_ keymem.key_mem\[3\]\[70\] _08009_ keymem.key_mem\[9\]\[70\]
+ _07705_ _08402_ sky130_fd_sc_hd__a221o_2
XFILLER_0_5_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_150_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14608_ VGND VPWR VGND VPWR _10075_ _10056_ keymem.round_ctr_reg\[0\] _10076_ sky130_fd_sc_hd__a21o_2
XFILLER_0_28_344 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18376_ VPWR VGND VGND VPWR _04270_ _04194_ _04268_ sky130_fd_sc_hd__nand2_2
X_15588_ _10215_ _11046_ keymem.prev_key1_reg\[110\] _10229_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_145_349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_44_826 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17327_ VPWR VGND VGND VPWR _02750_ _03420_ keymem.prev_key0_reg\[91\] sky130_fd_sc_hd__nor2_2
XFILLER_0_56_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14539_ VGND VPWR VGND VPWR _10007_ _09204_ _09211_ _09107_ _09658_ _10006_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_50_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_70_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17258_ VGND VPWR VGND VPWR _02461_ _02460_ _03358_ keymem.prev_key0_reg\[84\] sky130_fd_sc_hd__a21oi_2
XFILLER_0_148_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_153_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16209_ VPWR VGND VGND VPWR _11245_ _11238_ _02374_ _11372_ _11257_ sky130_fd_sc_hd__o22ai_2
X_17189_ VGND VPWR VPWR VGND _03296_ keymem.key_mem\[14\]\[76\] _03295_ _03297_ sky130_fd_sc_hd__mux2_2
XFILLER_0_113_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_767 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_109_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_256_913 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_227_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_242_106 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22910_ VGND VPWR VGND VPWR _02194_ _06911_ _06882_ keymem.prev_key1_reg\[17\] sky130_fd_sc_hd__o21a_2
XFILLER_0_166_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_38_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23890_ VGND VPWR VPWR VGND clk _00383_ reset_n keymem.key_mem\[13\]\[11\] sky130_fd_sc_hd__dfrtp_2
X_22841_ VPWR VGND VGND VPWR _06869_ keymem.rcon_reg\[3\] keymem.rcon_logic.tmp_rcon\[0\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_194_1191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_250_150 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_17_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25560_ VGND VPWR VPWR VGND clk _02053_ reset_n keymem.key_mem\[0\]\[17\] sky130_fd_sc_hd__dfrtp_2
X_22772_ VGND VPWR _02119_ _06848_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24511_ VGND VPWR VPWR VGND clk _01004_ reset_n keymem.key_mem\[9\]\[120\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_195_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_194_1_Right_795 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_93_203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21723_ VGND VPWR _01587_ _06331_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25491_ VGND VPWR VPWR VGND clk _01984_ reset_n keymem.key_mem\[1\]\[76\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24442_ VGND VPWR VPWR VGND clk _00935_ reset_n keymem.key_mem\[9\]\[51\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_344 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21654_ VGND VPWR VPWR VGND _06286_ _02861_ keymem.key_mem\[4\]\[31\] _06295_ sky130_fd_sc_hd__mux2_2
XFILLER_0_46_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20605_ VGND VPWR _05736_ _05679_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_35_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24373_ VGND VPWR VPWR VGND clk _00866_ reset_n keymem.key_mem\[10\]\[110\] sky130_fd_sc_hd__dfrtp_2
X_21585_ VGND VPWR VGND VPWR keymem.round_ctr_reg\[3\] _06257_ keymem.key_mem_we keymem.round_ctr_reg\[2\]
+ _08925_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_46_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_62_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23324_ VPWR VGND _07203_ _07128_ enc_block.block_w2_reg\[4\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_20536_ VGND VPWR VPWR VGND _05692_ _02479_ keymem.key_mem\[8\]\[20\] _05700_ sky130_fd_sc_hd__mux2_2
XFILLER_0_127_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23255_ VPWR VGND _07141_ enc_block.block_w3_reg\[29\] enc_block.block_w3_reg\[28\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_127_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20467_ VGND VPWR VPWR VGND _05660_ _03592_ keymem.key_mem\[9\]\[116\] _05663_ sky130_fd_sc_hd__mux2_2
XFILLER_0_28_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22206_ VGND VPWR _01811_ _06590_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_162_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_762 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23186_ VGND VPWR VGND VPWR _03650_ _03649_ _03653_ _07080_ sky130_fd_sc_hd__a21o_2
XFILLER_0_28_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20398_ VGND VPWR _00967_ _05626_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22137_ VGND VPWR _06553_ _06552_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_203_1154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_98_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_467 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22068_ VGND VPWR _06516_ _06402_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_238_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13910_ VPWR VGND VPWR VGND _09299_ _09317_ _09300_ _09297_ _09382_ sky130_fd_sc_hd__or4_2
X_21019_ VGND VPWR VPWR VGND _05956_ _05069_ keymem.key_mem\[7\]\[117\] _05958_ sky130_fd_sc_hd__mux2_2
X_14890_ VGND VPWR VGND VPWR _09646_ _09127_ _09124_ _09204_ _10355_ sky130_fd_sc_hd__o22a_2
X_13841_ VGND VPWR VGND VPWR _09305_ _09302_ _09313_ _09312_ sky130_fd_sc_hd__a21oi_2
X_25827_ VGND VPWR VPWR VGND clk _02320_ reset_n enc_block.block_w3_reg\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_199_555 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_138_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_134_1215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_35_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13772_ VPWR VGND VPWR VGND _09244_ enc_block.block_w0_reg\[24\] _08995_ sky130_fd_sc_hd__or2_2
XFILLER_0_39_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16560_ VGND VPWR VPWR VGND _02719_ _02708_ _02715_ _02716_ _02718_ sky130_fd_sc_hd__o31a_2
X_25758_ keymem.prev_key1_reg\[74\] clk _02251_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_35_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15511_ VPWR VGND VGND VPWR _10971_ key[140] _10091_ sky130_fd_sc_hd__nand2_2
X_24709_ VGND VPWR VPWR VGND clk _01202_ reset_n keymem.key_mem\[7\]\[62\] sky130_fd_sc_hd__dfrtp_2
X_12723_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[56\] _07919_ keymem.key_mem\[8\]\[56\]
+ _08211_ _08270_ sky130_fd_sc_hd__a22o_2
X_16491_ VGND VPWR VGND VPWR _11141_ _11113_ keymem.prev_key1_reg\[119\] _02652_ sky130_fd_sc_hd__a21o_2
X_25689_ keymem.prev_key1_reg\[5\] clk _02182_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_18230_ VPWR VGND VGND VPWR _04137_ _04004_ _11142_ sky130_fd_sc_hd__nand2_2
X_15442_ VGND VPWR VGND VPWR _09981_ _09941_ keymem.prev_key1_reg\[107\] _10903_ sky130_fd_sc_hd__a21o_2
X_12654_ VPWR VGND VPWR VGND _08207_ keymem.key_mem\[6\]\[49\] _07711_ keymem.key_mem\[9\]\[49\]
+ _07705_ _08208_ sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_68_1_Right_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_242_77 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_84_269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_127_349 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18161_ VGND VPWR VPWR VGND _03974_ enc_block.block_w0_reg\[8\] _04074_ _04075_ sky130_fd_sc_hd__mux2_2
X_12585_ VGND VPWR _08145_ _07534_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15373_ VPWR VGND VPWR VGND _10834_ _10826_ _10825_ key[138] _09544_ _10835_ sky130_fd_sc_hd__a221o_2
XFILLER_0_154_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17112_ VPWR VGND VGND VPWR _03228_ keymem.key_mem\[14\]\[68\] _09541_ sky130_fd_sc_hd__nand2_2
X_14324_ VGND VPWR VPWR VGND _09793_ _09731_ _09728_ _09794_ sky130_fd_sc_hd__mux2_2
X_18092_ VGND VPWR _04011_ enc_block.block_w1_reg\[19\] enc_block.block_w0_reg\[27\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_145_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_149_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14255_ VGND VPWR VPWR VGND _09541_ keymem.key_mem\[14\]\[1\] _09725_ _09726_ sky130_fd_sc_hd__mux2_2
X_17043_ _02822_ _03165_ _02817_ _02824_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_12_Left_280 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_46_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13206_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[104\] _07610_ keymem.key_mem\[2\]\[104\]
+ _07547_ _08705_ sky130_fd_sc_hd__a22o_2
X_14186_ VGND VPWR VGND VPWR _09148_ _09216_ _09657_ _09069_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_106_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_586 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13137_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[97\] _07685_ keymem.key_mem\[4\]\[97\]
+ _07636_ _08643_ sky130_fd_sc_hd__a22o_2
X_18994_ VPWR VGND VPWR VGND _04825_ _04605_ _04823_ sky130_fd_sc_hd__or2_2
XFILLER_0_267_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13068_ VGND VPWR VGND VPWR _07835_ keymem.key_mem\[13\]\[90\] _08578_ _08580_ _08581_
+ _08480_ sky130_fd_sc_hd__a2111o_2
X_17945_ VGND VPWR _00246_ _03894_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_253_949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12019_ VGND VPWR _07621_ _07620_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17876_ VGND VPWR _00224_ _03847_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_79_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19615_ VGND VPWR _00600_ _05210_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_156_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16827_ VGND VPWR VPWR VGND _08927_ _02968_ key[170] _02969_ sky130_fd_sc_hd__mux2_2
XFILLER_0_233_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19546_ VGND VPWR VGND VPWR _05174_ keymem.key_mem_we _03217_ _05164_ _00567_ sky130_fd_sc_hd__a31o_2
XFILLER_0_57_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_215_1047 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16758_ VPWR VGND VGND VPWR _09988_ _02906_ key[36] sky130_fd_sc_hd__nor2_2
XFILLER_0_48_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_117_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15709_ VPWR VGND VPWR VGND _11165_ enc_block.block_w0_reg\[18\] _09273_ sky130_fd_sc_hd__or2_2
X_19477_ VGND VPWR VGND VPWR _05137_ keymem.key_mem_we _02904_ _05135_ _00535_ sky130_fd_sc_hd__a31o_2
X_16689_ VGND VPWR VPWR VGND _02620_ _02636_ _02613_ _02842_ sky130_fd_sc_hd__or3_2
XFILLER_0_14_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18428_ VGND VPWR VGND VPWR _04315_ _03992_ _04312_ _04313_ _00308_ sky130_fd_sc_hd__a31o_2
XFILLER_0_115_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18359_ VPWR VGND _04255_ _04254_ enc_block.round_key\[122\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_267_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_44_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21370_ VGND VPWR VPWR VGND _06140_ _02720_ keymem.key_mem\[5\]\[25\] _06145_ sky130_fd_sc_hd__mux2_2
XFILLER_0_185_1168 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_44_689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_128_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20321_ VGND VPWR _00930_ _05586_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_4_775 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_64_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23040_ VGND VPWR VPWR VGND _06960_ _06990_ keymem.prev_key1_reg\[68\] _06991_ sky130_fd_sc_hd__mux2_2
X_20252_ VGND VPWR _00897_ _05550_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_25_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_101_249 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_204_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20183_ VGND VPWR VPWR VGND _05504_ _03560_ keymem.key_mem\[10\]\[111\] _05512_ sky130_fd_sc_hd__mux2_2
XFILLER_0_204_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24991_ VGND VPWR VPWR VGND clk _01484_ reset_n keymem.key_mem\[5\]\[88\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_239_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1264 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23942_ VGND VPWR VPWR VGND clk _00435_ reset_n keymem.key_mem\[13\]\[63\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_208_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23873_ VGND VPWR VPWR VGND clk _00366_ reset_n enc_block.block_w2_reg\[26\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_135_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25612_ VGND VPWR VPWR VGND clk _02105_ reset_n keymem.key_mem\[0\]\[69\] sky130_fd_sc_hd__dfrtp_2
X_22824_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[123\] _06839_ _03864_ _05081_ _02159_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_211_323 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_196_536 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_227 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_1029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22755_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[72\] _06837_ _06836_ _04986_ _02108_
+ sky130_fd_sc_hd__a22o_2
X_25543_ VGND VPWR VPWR VGND clk _02036_ reset_n keymem.key_mem\[0\]\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_439 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_215_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_211_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_195_1_Right_796 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21706_ VGND VPWR _01579_ _06322_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25474_ VGND VPWR VPWR VGND clk _01967_ reset_n keymem.key_mem\[1\]\[59\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22686_ VGND VPWR VPWR VGND _06809_ keymem.key_mem\[0\]\[31\] _02862_ _06815_ sky130_fd_sc_hd__mux2_2
XFILLER_0_109_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24425_ VGND VPWR VPWR VGND clk _00918_ reset_n keymem.key_mem\[9\]\[34\] sky130_fd_sc_hd__dfrtp_2
X_21637_ VGND VPWR _06286_ _06262_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_30_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24356_ VGND VPWR VPWR VGND clk _00849_ reset_n keymem.key_mem\[10\]\[93\] sky130_fd_sc_hd__dfrtp_2
X_12370_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[23\] _07587_ keymem.key_mem\[6\]\[23\]
+ _07771_ _07950_ sky130_fd_sc_hd__a22o_2
XFILLER_0_30_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21568_ VGND VPWR _01515_ _06248_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_117_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_34_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23307_ VPWR VGND VGND VPWR _07188_ _07185_ _07186_ sky130_fd_sc_hd__nand2_2
XFILLER_0_16_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_126_1_Left_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20519_ VGND VPWR VPWR VGND _05680_ _10976_ keymem.key_mem\[8\]\[12\] _05691_ sky130_fd_sc_hd__mux2_2
X_24287_ VGND VPWR VPWR VGND clk _00780_ reset_n keymem.key_mem\[10\]\[24\] sky130_fd_sc_hd__dfrtp_2
X_21499_ VGND VPWR _01482_ _06212_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14040_ VPWR VGND VGND VPWR _09511_ _09512_ _07378_ sky130_fd_sc_hd__nor2_2
X_23238_ VGND VPWR _07126_ _07092_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_30_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_570 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_222_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_372 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23169_ VGND VPWR _02295_ _07069_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_247_743 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_219_434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_776 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_140_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15991_ VGND VPWR _11447_ _11446_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_101_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_228_990 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17730_ VGND VPWR VPWR VGND _03723_ _02869_ keymem.prev_key0_reg\[32\] _03753_ sky130_fd_sc_hd__mux2_2
X_14942_ VGND VPWR VGND VPWR enc_block.block_w2_reg\[11\] _09269_ _10387_ _10404_
+ _10406_ _10405_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_261_234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_175_1348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17661_ VGND VPWR VPWR VGND _03703_ _03702_ keymem.prev_key0_reg\[12\] _03704_ sky130_fd_sc_hd__mux2_2
X_14873_ VGND VPWR VGND VPWR _09217_ _09077_ _09102_ _09099_ _10338_ sky130_fd_sc_hd__o22a_2
XFILLER_0_215_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19400_ VPWR VGND keymem.key_mem\[12\]\[0\] _05096_ _05095_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16612_ VGND VPWR VGND VPWR keymem.rcon_logic.tmp_rcon\[5\] _02430_ _02768_ _02458_
+ sky130_fd_sc_hd__a21bo_2
X_13824_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[27\] _08969_ _09296_ _09251_ _08964_
+ _09252_ sky130_fd_sc_hd__a32oi_2
X_17592_ VPWR VGND VGND VPWR _03651_ _02801_ _02802_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19331_ VPWR VGND keymem.key_mem_we _05048_ _03538_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_159_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16543_ VPWR VGND VGND VPWR _02702_ _02696_ _02701_ sky130_fd_sc_hd__nand2_2
X_13755_ VPWR VGND VPWR VGND _09226_ _09227_ _09224_ _09225_ sky130_fd_sc_hd__or3b_2
XFILLER_0_6_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19262_ VPWR VGND keymem.key_mem\[13\]\[82\] _05004_ _04979_ VPWR VGND sky130_fd_sc_hd__and2_2
X_12706_ VGND VPWR VGND VPWR _08255_ _07958_ keymem.key_mem\[8\]\[54\] _08254_ _07746_
+ sky130_fd_sc_hd__a211o_2
X_16474_ VPWR VGND VGND VPWR _11414_ _02632_ _02633_ _02634_ _02635_ sky130_fd_sc_hd__and4b_2
X_13686_ VGND VPWR VGND VPWR _09156_ _09097_ _09138_ _09157_ _09158_ sky130_fd_sc_hd__o22a_2
XFILLER_0_57_269 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_461 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18213_ _04120_ _04122_ _04065_ _04121_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_186_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15425_ VGND VPWR VGND VPWR _10510_ _10449_ _10886_ _10507_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_112_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19193_ VGND VPWR VGND VPWR _04962_ keymem.key_mem_we _03091_ _04924_ _00426_ sky130_fd_sc_hd__a31o_2
X_12637_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[48\] _07919_ keymem.key_mem\[4\]\[48\]
+ _07693_ _08192_ sky130_fd_sc_hd__a22o_2
XFILLER_0_26_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_142_105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18144_ _04057_ _04059_ _04008_ _04058_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_245_1018 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_976 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15356_ VGND VPWR keymem.prev_key0_reg\[106\] _10815_ _10818_ _10816_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_12568_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[41\] _07760_ keymem.key_mem\[8\]\[41\]
+ _07878_ _08130_ sky130_fd_sc_hd__a22o_2
XFILLER_0_198_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_186_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_1173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14307_ VPWR VGND VGND VPWR _09565_ _09777_ _09268_ sky130_fd_sc_hd__nor2_2
X_18075_ VPWR VGND VPWR VGND _03995_ _03992_ _03991_ enc_block.block_w0_reg\[1\] _03976_
+ _00275_ sky130_fd_sc_hd__a221o_2
X_15287_ VPWR VGND VPWR VGND _10749_ _10528_ _10508_ sky130_fd_sc_hd__or2_2
X_12499_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[35\] _07918_ keymem.key_mem\[11\]\[35\]
+ _07658_ _08067_ sky130_fd_sc_hd__a22o_2
X_17026_ VGND VPWR _03150_ _03149_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_145_1163 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_22_862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14238_ VGND VPWR VGND VPWR _09708_ _09679_ _07386_ _09709_ sky130_fd_sc_hd__a21o_2
XFILLER_0_21_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14169_ VPWR VGND VGND VPWR _09145_ _09121_ _09640_ _09173_ _09081_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_42_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18977_ VGND VPWR _04810_ _04808_ _04809_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_237_275 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_256_1114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_252_212 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_56_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17928_ VGND VPWR VGND VPWR _03489_ keymem.prev_key1_reg\[100\] _03883_ _03818_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_253_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_256_1158 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_193_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17859_ VGND VPWR _03836_ _03673_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_234_1423 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20870_ VPWR VGND keymem.key_mem\[7\]\[47\] _05879_ _05856_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_95_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_191_1172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_152_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19529_ VGND VPWR VGND VPWR _05165_ keymem.key_mem_we _03140_ _05164_ _00559_ sky130_fd_sc_hd__a31o_2
XFILLER_0_88_394 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_18_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22540_ VGND VPWR _01977_ _06758_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_220_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_834 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_130_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_29_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_191_1_Left_458 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_867 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_612 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22471_ VGND VPWR VPWR VGND _06726_ keymem.key_mem\[1\]\[29\] _02812_ _06730_ sky130_fd_sc_hd__mux2_2
XFILLER_0_9_889 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_130_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24210_ VGND VPWR VPWR VGND clk _00703_ reset_n keymem.key_mem\[11\]\[75\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_8_388 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21422_ VGND VPWR VPWR VGND _06162_ _03056_ keymem.key_mem\[5\]\[50\] _06172_ sky130_fd_sc_hd__mux2_2
XFILLER_0_173_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25190_ VGND VPWR VPWR VGND clk _01683_ reset_n keymem.key_mem\[3\]\[31\] sky130_fd_sc_hd__dfrtp_2
X_24141_ VGND VPWR VPWR VGND clk _00634_ reset_n keymem.key_mem\[11\]\[6\] sky130_fd_sc_hd__dfrtp_2
X_21353_ VGND VPWR VPWR VGND _06128_ _11546_ keymem.key_mem\[5\]\[17\] _06136_ sky130_fd_sc_hd__mux2_2
XFILLER_0_31_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_572 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20304_ VGND VPWR _00922_ _05577_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24072_ VGND VPWR VPWR VGND clk _00565_ reset_n keymem.key_mem\[12\]\[65\] sky130_fd_sc_hd__dfrtp_2
X_21284_ VGND VPWR _06098_ _05970_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_141_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23023_ VPWR VGND VGND VPWR _06981_ _03156_ _06976_ sky130_fd_sc_hd__nand2_2
X_20235_ VGND VPWR _00889_ _05541_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_97_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_99_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_905 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_1257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_204_1282 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_228_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20166_ VGND VPWR VPWR VGND _05493_ _03511_ keymem.key_mem\[10\]\[103\] _05503_ sky130_fd_sc_hd__mux2_2
XFILLER_0_141_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_244_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_196_1061 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24974_ VGND VPWR VPWR VGND clk _01467_ reset_n keymem.key_mem\[5\]\[71\] sky130_fd_sc_hd__dfrtp_2
X_20097_ VGND VPWR VPWR VGND _05457_ _03245_ keymem.key_mem\[10\]\[70\] _05467_ sky130_fd_sc_hd__mux2_2
X_23925_ VGND VPWR VPWR VGND clk _00418_ reset_n keymem.key_mem\[13\]\[46\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_224_470 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_58_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11870_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[6\] dec_new_block\[102\]
+ _07499_ sky130_fd_sc_hd__mux2_2
X_23856_ VGND VPWR VPWR VGND clk _00349_ reset_n enc_block.block_w2_reg\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22807_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[108\] _06858_ _06857_ _05050_ _02144_
+ sky130_fd_sc_hd__a22o_2
X_23787_ VGND VPWR VPWR VGND clk _00280_ reset_n enc_block.block_w0_reg\[6\] sky130_fd_sc_hd__dfrtp_2
X_20999_ VGND VPWR _01247_ _05947_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_39_258 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13540_ VPWR VGND VGND VPWR _09011_ _09012_ _09007_ sky130_fd_sc_hd__nor2_2
XFILLER_0_109_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25526_ VGND VPWR VPWR VGND clk _02019_ reset_n keymem.key_mem\[1\]\[111\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_109_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22738_ VGND VPWR _02099_ _06834_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_55_729 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13471_ VGND VPWR _08943_ _08942_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_109_146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25457_ VGND VPWR VPWR VGND clk _01950_ reset_n keymem.key_mem\[1\]\[42\] sky130_fd_sc_hd__dfrtp_2
X_22669_ VGND VPWR VPWR VGND _06798_ keymem.key_mem\[0\]\[23\] _02661_ _06806_ sky130_fd_sc_hd__mux2_2
X_15210_ VPWR VGND VGND VPWR _10646_ _10672_ _10673_ _10588_ _10568_ _10535_ sky130_fd_sc_hd__o32ai_2
X_12422_ VGND VPWR VGND VPWR _07924_ keymem.key_mem\[9\]\[28\] _07994_ _07996_ _07997_
+ _07662_ sky130_fd_sc_hd__a2111o_2
X_24408_ VGND VPWR VPWR VGND clk _00901_ reset_n keymem.key_mem\[9\]\[17\] sky130_fd_sc_hd__dfrtp_2
X_16190_ VPWR VGND VPWR VGND _02352_ _02354_ _02355_ _11616_ _02351_ sky130_fd_sc_hd__or4b_2
XFILLER_0_1_1460 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25388_ VGND VPWR VPWR VGND clk _01881_ reset_n keymem.key_mem\[2\]\[101\] sky130_fd_sc_hd__dfrtp_2
X_15141_ VPWR VGND VGND VPWR _10595_ _10602_ _10605_ _10489_ _10604_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_62_272 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12353_ VGND VPWR enc_block.round_key\[21\] _07934_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_129_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24339_ VGND VPWR VPWR VGND clk _00832_ reset_n keymem.key_mem\[10\]\[76\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_132_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15072_ VGND VPWR _10536_ _10535_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_105_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_107_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12284_ VGND VPWR enc_block.round_key\[16\] _07870_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_10_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14023_ VGND VPWR _09495_ _09400_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18900_ VGND VPWR VGND VPWR _04740_ _04505_ _04738_ _04739_ _04741_ sky130_fd_sc_hd__a31o_2
XFILLER_0_120_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19880_ VGND VPWR _00724_ _05351_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_205_1079 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18831_ VPWR VGND VPWR VGND _04678_ block[40] _03980_ enc_block.block_w0_reg\[8\]
+ _03978_ _04679_ sky130_fd_sc_hd__a221o_2
XFILLER_0_248_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18762_ VGND VPWR _04616_ enc_block.block_w2_reg\[25\] enc_block.block_w0_reg\[10\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15974_ _11287_ _11430_ _11356_ _11408_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_179_1292 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_218_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1145 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17713_ VPWR VGND VGND VPWR _03741_ _03742_ _03731_ sky130_fd_sc_hd__nor2_2
X_14925_ VGND VPWR VGND VPWR _10389_ enc_block.sword_ctr_reg\[0\] enc_block.block_w1_reg\[9\]
+ enc_block.sword_ctr_reg\[1\] sky130_fd_sc_hd__and3b_2
X_18693_ VPWR VGND VGND VPWR _04554_ _04341_ _04553_ sky130_fd_sc_hd__nand2_2
XFILLER_0_264_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1226 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_76_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17644_ VGND VPWR VPWR VGND _03691_ key[135] keymem.prev_key1_reg\[7\] _03692_ sky130_fd_sc_hd__mux2_2
XFILLER_0_264_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14856_ VGND VPWR VGND VPWR _10318_ _10287_ _10320_ _10321_ sky130_fd_sc_hd__a21o_2
XFILLER_0_118_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13807_ VPWR VGND VPWR VGND _09279_ enc_block.block_w0_reg\[30\] _08952_ sky130_fd_sc_hd__or2_2
XFILLER_0_202_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17575_ VGND VPWR VGND VPWR _03636_ _02928_ _02877_ key[123] sky130_fd_sc_hd__o21a_2
XFILLER_0_15_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14787_ VGND VPWR VGND VPWR _09343_ _09366_ _09335_ _09403_ _10253_ sky130_fd_sc_hd__o22a_2
X_11999_ VGND VPWR _07602_ _07601_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19314_ VGND VPWR _00473_ _05036_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16526_ VPWR VGND VPWR VGND _02686_ key[152] _10286_ sky130_fd_sc_hd__or2_2
X_13738_ VPWR VGND VPWR VGND _09044_ _08997_ _09034_ _08977_ _09210_ sky130_fd_sc_hd__or4_2
XFILLER_0_133_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19245_ VGND VPWR _04993_ _04876_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16457_ VPWR VGND VGND VPWR _11385_ _02618_ _11257_ sky130_fd_sc_hd__nor2_2
X_13669_ VGND VPWR _09141_ _09050_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_229_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15408_ VPWR VGND VGND VPWR _10868_ _10869_ _10866_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19176_ VGND VPWR VPWR VGND _04951_ _04950_ keymem.key_mem\[13\]\[48\] _04952_ sky130_fd_sc_hd__mux2_2
XFILLER_0_170_211 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_60_209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16388_ VGND VPWR VPWR VGND _11041_ keymem.key_mem\[14\]\[21\] _02550_ _02551_ sky130_fd_sc_hd__mux2_2
XFILLER_0_229_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18127_ VPWR VGND VPWR VGND _04043_ _04040_ _04039_ enc_block.block_w0_reg\[5\] _03976_
+ _00279_ sky130_fd_sc_hd__a221o_2
X_15339_ VGND VPWR VGND VPWR _10800_ _10799_ _10801_ _10798_ _10796_ sky130_fd_sc_hd__nand4_2
XFILLER_0_53_294 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_83_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1282 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18058_ VGND VPWR _03979_ _03956_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_13_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_123_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17009_ VPWR VGND VPWR VGND _03134_ keymem.prev_key1_reg\[59\] sky130_fd_sc_hd__inv_2
XFILLER_0_10_832 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_201_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20020_ VGND VPWR VPWR VGND _05424_ _02883_ keymem.key_mem\[10\]\[33\] _05427_ sky130_fd_sc_hd__mux2_2
XFILLER_0_158_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_123_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_203_Right_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_94_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21971_ VGND VPWR VPWR VGND _06462_ _04955_ keymem.key_mem\[3\]\[50\] _06465_ sky130_fd_sc_hd__mux2_2
XFILLER_0_154_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23710_ keymem.prev_key0_reg\[66\] clk _00207_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20922_ VPWR VGND keymem.key_mem\[7\]\[71\] _05907_ _05899_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_94_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24690_ VGND VPWR VPWR VGND clk _01183_ reset_n keymem.key_mem\[7\]\[43\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_55_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_68_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_90_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20853_ VGND VPWR _01178_ _05870_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23641_ VGND VPWR VPWR VGND clk _00010_ reset_n keymem.key_mem_we sky130_fd_sc_hd__dfrtp_2
XFILLER_0_7_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23572_ VGND VPWR VPWR VGND clk _00073_ reset_n keymem.key_mem\[14\]\[61\] sky130_fd_sc_hd__dfrtp_2
X_20784_ VGND VPWR VPWR VGND _05820_ _04889_ keymem.key_mem\[7\]\[7\] _05833_ sky130_fd_sc_hd__mux2_2
XFILLER_0_193_358 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22523_ VGND VPWR VPWR VGND _06739_ keymem.key_mem\[1\]\[62\] _03173_ _06749_ sky130_fd_sc_hd__mux2_2
X_25311_ VGND VPWR VPWR VGND clk _01804_ reset_n keymem.key_mem\[2\]\[24\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_664 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_420 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_263 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_228_1002 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_212_Right_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25242_ VGND VPWR VPWR VGND clk _01735_ reset_n keymem.key_mem\[3\]\[83\] sky130_fd_sc_hd__dfrtp_2
X_22454_ VGND VPWR VPWR VGND _06715_ keymem.key_mem\[1\]\[21\] _02550_ _06721_ sky130_fd_sc_hd__mux2_2
XFILLER_0_146_285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_464 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_106_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21405_ VGND VPWR _01437_ _06163_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_165_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25173_ VGND VPWR VPWR VGND clk _01666_ reset_n keymem.key_mem\[3\]\[14\] sky130_fd_sc_hd__dfrtp_2
X_22385_ VGND VPWR VPWR VGND _06680_ _03600_ keymem.key_mem\[2\]\[117\] _06684_ sky130_fd_sc_hd__mux2_2
XFILLER_0_161_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_892 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24124_ VGND VPWR VPWR VGND clk _00617_ reset_n keymem.key_mem\[12\]\[117\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_607 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21336_ VGND VPWR VPWR VGND _06117_ _10746_ keymem.key_mem\[5\]\[9\] _06127_ sky130_fd_sc_hd__mux2_2
XFILLER_0_248_304 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_66_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24055_ VGND VPWR VPWR VGND clk _00548_ reset_n keymem.key_mem\[12\]\[48\] sky130_fd_sc_hd__dfrtp_2
X_21267_ VGND VPWR _01373_ _06089_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_60_1021 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_64_1190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23006_ VGND VPWR VPWR VGND _06960_ _03089_ keymem.prev_key1_reg\[54\] _06971_ sky130_fd_sc_hd__mux2_2
X_20218_ VPWR VGND VGND VPWR _05530_ keymem.key_mem_we keymem.round_ctr_reg\[0\] sky130_fd_sc_hd__nand2_2
XFILLER_0_102_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_263_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21198_ VGND VPWR _01340_ _06053_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_198_1167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_221_Right_90 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20149_ VGND VPWR _00850_ _05494_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_102_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24957_ VGND VPWR VPWR VGND clk _01450_ reset_n keymem.key_mem\[5\]\[54\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_235_1017 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12971_ VGND VPWR VGND VPWR _08494_ _07593_ keymem.key_mem\[9\]\[80\] _08491_ _08493_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_176_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14710_ VGND VPWR VGND VPWR _09216_ _09099_ _09089_ _09140_ _10177_ sky130_fd_sc_hd__o22a_2
XFILLER_0_73_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23908_ VGND VPWR VPWR VGND clk _00401_ reset_n keymem.key_mem\[13\]\[29\] sky130_fd_sc_hd__dfrtp_2
X_11922_ VGND VPWR VPWR VGND encdec enc_block.round\[0\] dec_round_nr\[0\] _07525_
+ sky130_fd_sc_hd__mux2_2
X_15690_ VGND VPWR VPWR VGND _09796_ key[15] _11147_ _11146_ _11145_ sky130_fd_sc_hd__o211a_2
X_24888_ VGND VPWR VPWR VGND clk _01381_ reset_n keymem.key_mem\[6\]\[113\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_169_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_197_653 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_73_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14641_ VPWR VGND VGND VPWR _09557_ _10069_ _10107_ _10108_ sky130_fd_sc_hd__nor3_2
X_11853_ VGND VPWR result[93] _07490_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23839_ VGND VPWR VPWR VGND clk _00332_ reset_n enc_block.block_w1_reg\[24\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_197_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17360_ VPWR VGND VGND VPWR _09732_ _03450_ key[222] sky130_fd_sc_hd__nor2_2
X_14572_ VGND VPWR VGND VPWR _09295_ _09248_ _10034_ _10039_ _10040_ _09345_ sky130_fd_sc_hd__a2111o_2
X_11784_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[27\] dec_new_block\[59\]
+ _07456_ sky130_fd_sc_hd__mux2_2
XFILLER_0_184_336 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_184_347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16311_ VPWR VGND VGND VPWR _02474_ _02475_ _02473_ sky130_fd_sc_hd__nor2_2
X_13523_ VGND VPWR _08995_ _08951_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_113_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25509_ VGND VPWR VPWR VGND clk _02002_ reset_n keymem.key_mem\[1\]\[94\] sky130_fd_sc_hd__dfrtp_2
X_17291_ VPWR VGND VGND VPWR _03388_ _02640_ _02641_ sky130_fd_sc_hd__nand2_2
XFILLER_0_32_1178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19030_ VPWR VGND VPWR VGND _04856_ _04103_ enc_block.block_w2_reg\[29\] _03952_
+ _04857_ sky130_fd_sc_hd__a22o_2
XFILLER_0_246_1102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16242_ VPWR VGND VGND VPWR _02403_ _02407_ _10092_ sky130_fd_sc_hd__nor2_2
XFILLER_0_42_209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_250_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13454_ VGND VPWR VPWR VGND keymem.round_ctr_reg\[3\] _08925_ keymem.round_ctr_reg\[2\]
+ _08926_ sky130_fd_sc_hd__or3_2
XFILLER_0_187_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12405_ VGND VPWR VGND VPWR _07982_ _07800_ keymem.key_mem\[1\]\[26\] _07979_ _07981_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_207_1108 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_183_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_829 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13385_ VGND VPWR enc_block.round_key\[121\] _08866_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16173_ VPWR VGND VPWR VGND _02338_ _09638_ _11559_ key[146] _11043_ _02339_ sky130_fd_sc_hd__a221o_2
XFILLER_0_84_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15124_ VGND VPWR _10588_ _10587_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_23_467 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_50_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_50_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12336_ VGND VPWR _07919_ _07918_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_80_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15055_ VGND VPWR _10519_ _10518_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_120_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_267_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12267_ VGND VPWR _07855_ _07556_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19932_ VGND VPWR _00749_ _05378_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14006_ VPWR VGND VGND VPWR _09362_ _09478_ _09447_ sky130_fd_sc_hd__nor2_2
X_19863_ VGND VPWR _00716_ _05342_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12198_ VGND VPWR VGND VPWR _07791_ _07650_ keymem.key_mem\[7\]\[10\] _07790_ _07572_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_120_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18814_ VGND VPWR _04664_ _03949_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19794_ VGND VPWR _00683_ _05306_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_120_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1242 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_21_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_194_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18745_ VGND VPWR VPWR VGND _04600_ enc_block.block_w2_reg\[0\] _03971_ _04601_ sky130_fd_sc_hd__mux2_2
X_15957_ _11412_ _11413_ _11266_ _11390_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_222_204 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_190_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_155_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_204_941 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_91_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_144_12 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14908_ VPWR VGND _10372_ keymem.prev_key1_reg\[40\] keymem.prev_key1_reg\[8\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
X_18676_ VPWR VGND VGND VPWR _04538_ _04539_ _04478_ sky130_fd_sc_hd__nor2_2
X_15888_ VGND VPWR _11344_ _11343_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_37_1034 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_91_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17627_ VGND VPWR VPWR VGND _03679_ key[130] keymem.prev_key1_reg\[2\] _03680_ sky130_fd_sc_hd__mux2_2
X_14839_ VPWR VGND VGND VPWR _09415_ _10304_ _09754_ sky130_fd_sc_hd__nor2_2
XFILLER_0_231_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17558_ VGND VPWR _00132_ _03621_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_19_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_175_358 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16509_ _11301_ _02669_ keymem.rcon_reg\[0\] _11438_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_131_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17489_ VGND VPWR _00123_ _03561_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19228_ VGND VPWR VGND VPWR _04982_ keymem.key_mem_we _03235_ _04968_ _00441_ sky130_fd_sc_hd__a31o_2
XPHY_EDGE_ROW_4_Left_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_913 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19159_ VGND VPWR _00414_ _04940_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_456 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22170_ VGND VPWR _01794_ _06571_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_242_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21121_ VGND VPWR VPWR VGND _06007_ _02913_ keymem.key_mem\[6\]\[36\] _06013_ sky130_fd_sc_hd__mux2_2
XFILLER_0_68_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_258_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1_383 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_159_1_Right_760 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21052_ VGND VPWR _01271_ _05976_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_266_690 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20003_ VGND VPWR VPWR VGND _05413_ _02721_ keymem.key_mem\[10\]\[25\] _05418_ sky130_fd_sc_hd__mux2_2
X_24811_ VGND VPWR VPWR VGND clk _01304_ reset_n keymem.key_mem\[6\]\[36\] sky130_fd_sc_hd__dfrtp_2
X_25791_ keymem.prev_key1_reg\[107\] clk _02284_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_20_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_59_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24742_ VGND VPWR VPWR VGND clk _01235_ reset_n keymem.key_mem\[7\]\[95\] sky130_fd_sc_hd__dfrtp_2
X_21954_ VGND VPWR VPWR VGND _06449_ _04939_ keymem.key_mem\[3\]\[42\] _06456_ sky130_fd_sc_hd__mux2_2
XFILLER_0_213_259 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_94_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20905_ VPWR VGND keymem.key_mem\[7\]\[63\] _05898_ _05886_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_178_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24673_ VGND VPWR VPWR VGND clk _01166_ reset_n keymem.key_mem\[7\]\[26\] sky130_fd_sc_hd__dfrtp_2
X_21885_ VGND VPWR VGND VPWR _06418_ keymem.key_mem_we _10836_ _06404_ _01662_ sky130_fd_sc_hd__a31o_2
XFILLER_0_16_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_103_2_Left_574 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_221_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20836_ VPWR VGND keymem.key_mem\[7\]\[31\] _05861_ _05856_ VPWR VGND sky130_fd_sc_hd__and2_2
X_23624_ VGND VPWR VPWR VGND clk _00125_ reset_n keymem.key_mem\[14\]\[113\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_64_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_49_386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_537 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23555_ VGND VPWR VPWR VGND clk _00056_ reset_n keymem.key_mem\[14\]\[44\] sky130_fd_sc_hd__dfrtp_2
X_20767_ VGND VPWR _05823_ _05822_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_18_751 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22506_ VGND VPWR VPWR VGND _06739_ keymem.key_mem\[1\]\[53\] _03083_ _06741_ sky130_fd_sc_hd__mux2_2
XFILLER_0_24_209 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23486_ VPWR VGND _07348_ _07347_ enc_block.round_key\[29\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_91_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20698_ VGND VPWR VPWR VGND _05783_ _03474_ keymem.key_mem\[8\]\[97\] _05785_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_220_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25225_ VGND VPWR VPWR VGND clk _01718_ reset_n keymem.key_mem\[3\]\[66\] sky130_fd_sc_hd__dfrtp_2
X_22437_ VGND VPWR VPWR VGND _06702_ keymem.key_mem\[1\]\[13\] _11040_ _06712_ sky130_fd_sc_hd__mux2_2
XFILLER_0_134_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_231 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_32_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13170_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[100\] _07593_ keymem.key_mem\[11\]\[100\]
+ _07838_ _08673_ sky130_fd_sc_hd__a22o_2
XFILLER_0_27_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25156_ VGND VPWR VPWR VGND clk _01649_ reset_n keymem.key_mem\[4\]\[125\] sky130_fd_sc_hd__dfrtp_2
X_22368_ VGND VPWR VPWR VGND _06669_ _03550_ keymem.key_mem\[2\]\[109\] _06675_ sky130_fd_sc_hd__mux2_2
XFILLER_0_20_415 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12121_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[6\] _07649_ keymem.key_mem\[11\]\[6\]
+ _07658_ _07718_ sky130_fd_sc_hd__a22o_2
X_24107_ VGND VPWR VPWR VGND clk _00600_ reset_n keymem.key_mem\[12\]\[100\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_206_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21319_ VGND VPWR _01396_ _06118_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_27_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25087_ VGND VPWR VPWR VGND clk _01580_ reset_n keymem.key_mem\[4\]\[56\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_202_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22299_ VGND VPWR VPWR VGND _06634_ _03295_ keymem.key_mem\[2\]\[76\] _06639_ sky130_fd_sc_hd__mux2_2
XFILLER_0_102_174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12052_ VGND VPWR _07652_ _07651_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24038_ VGND VPWR VPWR VGND clk _00531_ reset_n keymem.key_mem\[12\]\[31\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_229_381 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_263_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16860_ VGND VPWR _00056_ _02999_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_219_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15811_ VPWR VGND VPWR VGND _11266_ _11258_ _11180_ _11263_ _11267_ sky130_fd_sc_hd__or4_2
XFILLER_0_102_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_822 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_232_524 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16791_ VGND VPWR VPWR VGND _10363_ _10364_ _09516_ _02936_ sky130_fd_sc_hd__or3_2
XFILLER_0_99_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18530_ VPWR VGND _04408_ enc_block.block_w0_reg\[1\] enc_block.block_w2_reg\[18\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_137_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15742_ enc_block.sword_ctr_reg\[1\] _11198_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[21\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_12954_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[79\] _07649_ keymem.key_mem\[4\]\[79\]
+ _07636_ _08478_ sky130_fd_sc_hd__a22o_2
XFILLER_0_73_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_579 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_99_275 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_137_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11905_ VGND VPWR result[119] _07516_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18461_ VPWR VGND VGND VPWR _04346_ _04341_ _04344_ sky130_fd_sc_hd__nand2_2
X_15673_ VGND VPWR VGND VPWR _10628_ _10569_ _10627_ _10511_ _11130_ sky130_fd_sc_hd__o22a_2
XFILLER_0_197_461 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_73_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12885_ VGND VPWR VGND VPWR _07839_ keymem.key_mem\[11\]\[72\] _08413_ _08415_ _08416_
+ _07896_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_169_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_157_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_34_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17412_ VGND VPWR _03494_ key[101] _03495_ _03240_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_14624_ VGND VPWR _10092_ _10091_ VPWR VGND sky130_fd_sc_hd__buf_1
X_11836_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[21\] dec_new_block\[85\]
+ _07482_ sky130_fd_sc_hd__mux2_2
X_18392_ VPWR VGND VPWR VGND _04284_ _04189_ _04282_ enc_block.block_w0_reg\[29\]
+ _03993_ _00303_ sky130_fd_sc_hd__a221o_2
XFILLER_0_200_443 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_358 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17343_ VGND VPWR _03435_ _03434_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14555_ VPWR VGND VGND VPWR _09168_ _10023_ _09684_ sky130_fd_sc_hd__nor2_2
X_11767_ VGND VPWR result[50] _07447_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_200_498 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13506_ VPWR VGND VGND VPWR enc_block.block_w1_reg\[6\] enc_block.sword_ctr_reg\[0\]
+ _08978_ sky130_fd_sc_hd__or2b_2
XFILLER_0_99_17 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17274_ VGND VPWR VGND VPWR _03372_ _03371_ _03373_ keylen sky130_fd_sc_hd__a21oi_2
X_14486_ VPWR VGND VGND VPWR _09029_ _09147_ _09955_ _09124_ _09099_ sky130_fd_sc_hd__o22ai_2
X_11698_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[16\] dec_new_block\[16\]
+ _07413_ sky130_fd_sc_hd__mux2_2
XFILLER_0_148_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19013_ _04840_ _04842_ _04103_ _04841_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_16225_ VGND VPWR VGND VPWR _11250_ _11527_ _11336_ _11386_ _02390_ sky130_fd_sc_hd__o22a_2
XFILLER_0_125_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13437_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[127\] _07872_ keymem.key_mem\[8\]\[127\]
+ _07654_ _08913_ sky130_fd_sc_hd__a22o_2
XFILLER_0_10_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_905 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_140_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16156_ VGND VPWR VGND VPWR _11609_ _11395_ _11291_ _11426_ _11610_ sky130_fd_sc_hd__a31o_2
XFILLER_0_84_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_573 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_109_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13368_ VPWR VGND VPWR VGND _08850_ keymem.key_mem\[8\]\[120\] _08211_ keymem.key_mem\[4\]\[120\]
+ _07637_ _08851_ sky130_fd_sc_hd__a221o_2
XFILLER_0_140_247 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_23_286 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_267_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15107_ VGND VPWR VGND VPWR _10571_ _10564_ _10562_ _10567_ _10570_ sky130_fd_sc_hd__a211o_2
XFILLER_0_80_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12319_ VGND VPWR _07903_ _07539_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_45_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16087_ VGND VPWR VGND VPWR _09717_ _11540_ _11538_ _11539_ _11542_ sky130_fd_sc_hd__a31o_2
XFILLER_0_228_808 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13299_ VGND VPWR VGND VPWR _07648_ keymem.key_mem\[2\]\[113\] _08786_ _08788_ _08789_
+ _08736_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_224_1296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15038_ VPWR VGND VPWR VGND _10473_ _10409_ _10453_ _10451_ _10502_ sky130_fd_sc_hd__or4_2
X_19915_ VGND VPWR _00741_ _05369_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_267_498 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_48_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19846_ VGND VPWR _00708_ _05333_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_120_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_251_822 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19777_ VGND VPWR _00675_ _05297_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_263_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16989_ VPWR VGND VPWR VGND _03116_ key[185] _10322_ sky130_fd_sc_hd__or2_2
XFILLER_0_64_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_223_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_155_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18728_ VPWR VGND VGND VPWR _04585_ _04443_ _04584_ sky130_fd_sc_hd__nand2_2
XFILLER_0_56_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_155_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18659_ VPWR VGND VGND VPWR _04524_ _04307_ _04522_ sky130_fd_sc_hd__nand2_2
XFILLER_0_8_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_52_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21670_ VGND VPWR _01562_ _06303_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_59_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20621_ VGND VPWR _01072_ _05744_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_175_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23340_ VPWR VGND VPWR VGND _07217_ block[13] _03957_ enc_block.block_w1_reg\[13\]
+ _03952_ _07218_ sky130_fd_sc_hd__a221o_2
XFILLER_0_188_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20552_ VGND VPWR _01039_ _05708_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23271_ VPWR VGND VGND VPWR _07126_ _07156_ _04052_ sky130_fd_sc_hd__nor2_2
XFILLER_0_15_743 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_225_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20483_ VGND VPWR VPWR VGND _05534_ _03647_ keymem.key_mem\[9\]\[124\] _05671_ sky130_fd_sc_hd__mux2_2
XFILLER_0_15_754 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_116_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22222_ VGND VPWR _01819_ _06598_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25010_ VGND VPWR VPWR VGND clk _01503_ reset_n keymem.key_mem\[5\]\[107\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_30_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_127_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22153_ VGND VPWR VPWR VGND _06554_ _10369_ keymem.key_mem\[2\]\[7\] _06562_ sky130_fd_sc_hd__mux2_2
XFILLER_0_24_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_465 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21104_ VGND VPWR VPWR VGND _05996_ _02786_ keymem.key_mem\[6\]\[28\] _06004_ sky130_fd_sc_hd__mux2_2
X_22084_ VGND VPWR _01755_ _06524_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_203_1369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_58_Left_326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_239_690 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21035_ VGND VPWR VPWR VGND _05956_ _05085_ keymem.key_mem\[7\]\[125\] _05966_ sky130_fd_sc_hd__mux2_2
XFILLER_0_199_1284 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_242_800 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25843_ VGND VPWR VPWR VGND clk _02336_ reset_n enc_block.block_w3_reg\[31\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_177_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_173_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25774_ keymem.prev_key1_reg\[90\] clk _02267_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22986_ VGND VPWR _03013_ _03008_ _06959_ _03010_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_74_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_214_1410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24725_ VGND VPWR VPWR VGND clk _01218_ reset_n keymem.key_mem\[7\]\[78\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_70_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21937_ VPWR VGND keymem.key_mem\[3\]\[34\] _06447_ _06439_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_253_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12670_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[51\] _07845_ keymem.key_mem\[9\]\[51\]
+ _07919_ _08222_ sky130_fd_sc_hd__a22o_2
X_24656_ VGND VPWR VPWR VGND clk _01149_ reset_n keymem.key_mem\[7\]\[9\] sky130_fd_sc_hd__dfrtp_2
X_21868_ VGND VPWR VGND VPWR _06409_ keymem.key_mem_we _09862_ _06404_ _01654_ sky130_fd_sc_hd__a31o_2
XFILLER_0_210_1329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23607_ VGND VPWR VPWR VGND clk _00108_ reset_n keymem.key_mem\[14\]\[96\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_210_796 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20819_ VPWR VGND keymem.key_mem\[7\]\[23\] _05852_ _05844_ VPWR VGND sky130_fd_sc_hd__and2_2
X_21799_ VGND VPWR VPWR VGND _06366_ _03492_ keymem.key_mem\[4\]\[100\] _06371_ sky130_fd_sc_hd__mux2_2
X_24587_ VGND VPWR VPWR VGND clk _01080_ reset_n keymem.key_mem\[8\]\[68\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_181_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14340_ VGND VPWR VGND VPWR _09810_ _09001_ _09045_ _09015_ _09047_ _09809_ sky130_fd_sc_hd__a41o_2
XFILLER_0_147_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23538_ VGND VPWR VPWR VGND clk _00039_ reset_n keymem.key_mem\[14\]\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_110_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Right_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_184_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14271_ VPWR VGND VGND VPWR _09564_ _09466_ _09411_ _09399_ _09741_ _09740_ sky130_fd_sc_hd__o221a_2
XFILLER_0_0_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23469_ VGND VPWR _07333_ enc_block.round_key\[27\] _07332_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_145_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16010_ VPWR VGND VPWR VGND _11265_ _11258_ _11180_ _11167_ _11465_ sky130_fd_sc_hd__or4_2
XFILLER_0_184_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_122_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25208_ VGND VPWR VPWR VGND clk _01701_ reset_n keymem.key_mem\[3\]\[49\] sky130_fd_sc_hd__dfrtp_2
X_13222_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[105\] _07724_ keymem.key_mem\[2\]\[105\]
+ _07646_ _08720_ sky130_fd_sc_hd__a22o_2
XFILLER_0_81_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1269 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_145_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_584 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13153_ VGND VPWR VGND VPWR _08658_ _07712_ keymem.key_mem\[6\]\[98\] _08655_ _08657_
+ sky130_fd_sc_hd__a211o_2
X_25139_ VGND VPWR VPWR VGND clk _01632_ reset_n keymem.key_mem\[4\]\[108\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_42_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12104_ VGND VPWR _07702_ _07567_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17961_ VGND VPWR _00251_ _03905_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13084_ VGND VPWR enc_block.round_key\[91\] _08595_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_221_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16912_ VGND VPWR VPWR VGND _02986_ keymem.key_mem\[14\]\[49\] _03046_ _03047_ sky130_fd_sc_hd__mux2_2
X_19700_ VPWR VGND VGND VPWR _05257_ keymem.key_mem\[11\]\[11\] _05243_ sky130_fd_sc_hd__nand2_2
X_12035_ VGND VPWR _07636_ _07549_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_40_1244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17892_ VGND VPWR _03858_ _03395_ _00229_ _03675_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_178_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_256_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16843_ VPWR VGND VPWR VGND _02984_ _02979_ _02981_ _02982_ _02983_ _02496_ sky130_fd_sc_hd__o311a_2
X_19631_ VGND VPWR VPWR VGND _05216_ _05050_ keymem.key_mem\[12\]\[108\] _05219_ sky130_fd_sc_hd__mux2_2
XFILLER_0_260_630 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19562_ VGND VPWR VPWR VGND _00575_ _05095_ _03286_ _08922_ _05182_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_191_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16774_ VGND VPWR VGND VPWR _02921_ _10366_ _10187_ _10146_ sky130_fd_sc_hd__and3b_2
XFILLER_0_215_1207 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13986_ VPWR VGND VGND VPWR _09294_ _09458_ _09332_ sky130_fd_sc_hd__nor2_2
XFILLER_0_189_258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18513_ VGND VPWR _04393_ enc_block.block_w3_reg\[15\] _04392_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_152_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15725_ VGND VPWR VPWR VGND _11174_ _11180_ _11167_ _11181_ sky130_fd_sc_hd__or3_2
X_19493_ VGND VPWR VPWR VGND _05138_ _04941_ keymem.key_mem\[12\]\[43\] _05146_ sky130_fd_sc_hd__mux2_2
XFILLER_0_232_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12937_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[77\] _08016_ keymem.key_mem\[9\]\[77\]
+ _07593_ _08463_ sky130_fd_sc_hd__a22o_2
XFILLER_0_9_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_125_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18444_ VGND VPWR _04330_ _03979_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15656_ VGND VPWR VGND VPWR _10671_ _11112_ _11113_ _10551_ _10987_ sky130_fd_sc_hd__nor4_2
XFILLER_0_232_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12868_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[70\] _08391_ keymem.key_mem\[4\]\[70\]
+ _07692_ _08401_ sky130_fd_sc_hd__a22o_2
XFILLER_0_157_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_29_835 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14607_ VGND VPWR VGND VPWR _10065_ _10074_ _10075_ _10060_ _10070_ sky130_fd_sc_hd__nor4_2
X_18375_ VPWR VGND VPWR VGND _04269_ _04194_ _04268_ sky130_fd_sc_hd__or2_2
X_11819_ VGND VPWR result[76] _07473_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_5_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15587_ VGND VPWR VGND VPWR _10229_ _10215_ _11045_ keymem.prev_key1_reg\[110\] sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_56_Right_56 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12799_ VPWR VGND VPWR VGND _08338_ keymem.key_mem\[5\]\[63\] _07725_ keymem.key_mem\[1\]\[63\]
+ _07558_ _08339_ sky130_fd_sc_hd__a221o_2
XFILLER_0_126_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17326_ VGND VPWR _00102_ _03419_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14538_ VGND VPWR VGND VPWR _09097_ _09222_ _09110_ _09127_ _10006_ sky130_fd_sc_hd__o22a_2
XFILLER_0_43_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_160_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17257_ VGND VPWR _00095_ _03357_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14469_ VPWR VGND VGND VPWR _09102_ _09938_ _09134_ sky130_fd_sc_hd__nor2_2
XFILLER_0_226_1325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16208_ VPWR VGND VPWR VGND _02373_ _11485_ _11489_ sky130_fd_sc_hd__or2_2
XFILLER_0_52_860 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_113_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_148_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17188_ VGND VPWR _03296_ _09863_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_70_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_735 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_84_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16139_ VGND VPWR VGND VPWR _11283_ _11219_ _11593_ _11205_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_3_489 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_267_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_779 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_219_Left_486 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_200_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_209_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_208_351 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_196_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19829_ VGND VPWR _00700_ _05324_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_208_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_224_855 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22840_ VGND VPWR VGND VPWR keymem.rcon_reg\[3\] _06862_ _06868_ _06863_ _02167_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_251_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_196_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22771_ VGND VPWR VPWR VGND _06833_ keymem.key_mem\[0\]\[83\] _03356_ _06848_ sky130_fd_sc_hd__mux2_2
XFILLER_0_56_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_228_Left_495 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24510_ VGND VPWR VPWR VGND clk _01003_ reset_n keymem.key_mem\[9\]\[119\] sky130_fd_sc_hd__dfrtp_2
X_21722_ VGND VPWR VPWR VGND _06330_ _03183_ keymem.key_mem\[4\]\[63\] _06331_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25490_ VGND VPWR VPWR VGND clk _01983_ reset_n keymem.key_mem\[1\]\[75\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_8_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24441_ VGND VPWR VPWR VGND clk _00934_ reset_n keymem.key_mem\[9\]\[50\] sky130_fd_sc_hd__dfrtp_2
X_21653_ VGND VPWR _01554_ _06294_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20604_ VGND VPWR _01064_ _05735_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_266_1138 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21584_ VGND VPWR _01523_ _06256_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24372_ VGND VPWR VPWR VGND clk _00865_ reset_n keymem.key_mem\[10\]\[109\] sky130_fd_sc_hd__dfrtp_2
X_23323_ VGND VPWR _07202_ _04107_ _02316_ _07096_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_46_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20535_ VGND VPWR _01031_ _05699_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_144_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_61_145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_127_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_573 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23254_ VGND VPWR _07140_ enc_block.block_w1_reg\[13\] enc_block.block_w0_reg\[21\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20466_ VGND VPWR _00999_ _05662_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_166_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_584 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22205_ VGND VPWR VPWR VGND _06589_ _02861_ keymem.key_mem\[2\]\[31\] _06590_ sky130_fd_sc_hd__mux2_2
XFILLER_0_259_752 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_203_1100 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23185_ VGND VPWR VGND VPWR _02301_ _07079_ _06888_ keymem.prev_key1_reg\[124\] sky130_fd_sc_hd__o21a_2
X_20397_ VGND VPWR VPWR VGND _05614_ _03356_ keymem.key_mem\[9\]\[83\] _05626_ sky130_fd_sc_hd__mux2_2
XFILLER_0_24_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22136_ VGND VPWR _06552_ _06551_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_98_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_424 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22067_ VGND VPWR VGND VPWR _06515_ keymem.key_mem_we _03460_ _06498_ _01747_ sky130_fd_sc_hd__a31o_2
XFILLER_0_238_1229 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21018_ VGND VPWR _01256_ _05957_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_199_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13840_ VGND VPWR _09312_ _09311_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25826_ VGND VPWR VPWR VGND clk _02319_ reset_n enc_block.block_w3_reg\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_214_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_138_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13771_ VGND VPWR VGND VPWR enc_block.block_w1_reg\[24\] _08985_ _09022_ _09241_
+ _09243_ _09242_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_74_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1276 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25757_ keymem.prev_key1_reg\[73\] clk _02250_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_35_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22969_ VPWR VGND VPWR VGND _06949_ keymem.prev_key1_reg\[39\] _06926_ sky130_fd_sc_hd__or2_2
XFILLER_0_39_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15510_ VGND VPWR _10970_ keymem.prev_key1_reg\[12\] keymem.prev_key1_reg\[44\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24708_ VGND VPWR VPWR VGND clk _01201_ reset_n keymem.key_mem\[7\]\[61\] sky130_fd_sc_hd__dfrtp_2
X_12722_ VGND VPWR enc_block.round_key\[55\] _08269_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16490_ VGND VPWR VGND VPWR _11141_ keymem.prev_key1_reg\[119\] _02651_ _11113_ sky130_fd_sc_hd__nand3_2
XFILLER_0_35_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25688_ keymem.prev_key1_reg\[4\] clk _02181_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_15441_ VGND VPWR _10902_ _10328_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12653_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[49\] _07761_ keymem.key_mem\[1\]\[49\]
+ _07855_ _08207_ sky130_fd_sc_hd__a22o_2
X_24639_ VGND VPWR VPWR VGND clk _01132_ reset_n keymem.key_mem\[8\]\[120\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_154_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18160_ VPWR VGND VGND VPWR _10653_ _04074_ _04073_ sky130_fd_sc_hd__nor2_2
X_15372_ VPWR VGND VPWR VGND _10834_ _10325_ _10829_ _10830_ _10833_ _10281_ sky130_fd_sc_hd__o311a_2
X_12584_ VGND VPWR enc_block.round_key\[42\] _08144_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17111_ VGND VPWR _03227_ _03226_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_154_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14323_ VPWR VGND VGND VPWR _09793_ _09732_ _09792_ sky130_fd_sc_hd__nand2_2
X_18091_ VGND VPWR _04010_ enc_block.block_w2_reg\[11\] _04009_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17042_ VGND VPWR VGND VPWR _02822_ _02817_ _03164_ _02824_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_145_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1093 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14254_ VGND VPWR _09725_ _09724_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_81_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13205_ VGND VPWR enc_block.round_key\[103\] _08704_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_145_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_938 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14185_ VPWR VGND VGND VPWR _09166_ _09096_ _09656_ _09126_ _09121_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_96_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_42_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_249_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13136_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[97\] _07779_ keymem.key_mem\[1\]\[97\]
+ _07901_ _08642_ sky130_fd_sc_hd__a22o_2
XFILLER_0_21_598 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18993_ VPWR VGND VGND VPWR _04824_ _04605_ _04823_ sky130_fd_sc_hd__nand2_2
XFILLER_0_267_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13067_ VPWR VGND VPWR VGND _08579_ keymem.key_mem\[6\]\[90\] _07739_ keymem.key_mem\[10\]\[90\]
+ _07865_ _08580_ sky130_fd_sc_hd__a221o_2
X_17944_ VGND VPWR VPWR VGND _03874_ _03893_ keymem.prev_key0_reg\[105\] _03894_ sky130_fd_sc_hd__mux2_2
XFILLER_0_267_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12018_ VGND VPWR _07620_ _07576_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_178_1165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17875_ VGND VPWR VPWR VGND _03836_ _03846_ keymem.prev_key0_reg\[83\] _03847_ sky130_fd_sc_hd__mux2_2
X_19614_ VGND VPWR VPWR VGND _05205_ _05033_ keymem.key_mem\[12\]\[100\] _05210_ sky130_fd_sc_hd__mux2_2
XFILLER_0_79_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16826_ VPWR VGND _02968_ keymem.prev_key1_reg\[74\] keymem.prev_key1_reg\[42\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_117_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1332 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_156_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1015 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_92_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19545_ VPWR VGND keymem.key_mem\[12\]\[67\] _05174_ _05173_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_254_1086 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16757_ VGND VPWR _00047_ _02905_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13969_ VGND VPWR _09441_ _09440_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_117_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1059 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15708_ VGND VPWR VGND VPWR enc_block.block_w1_reg\[18\] _08947_ _10387_ _11162_
+ _11164_ _11163_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_243_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16688_ VPWR VGND VPWR VGND _11610_ _02611_ _02417_ _11481_ _02841_ sky130_fd_sc_hd__or4_2
XFILLER_0_53_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19476_ VPWR VGND keymem.key_mem\[12\]\[35\] _05137_ _05128_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_18_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18427_ VGND VPWR VPWR VGND _04314_ enc_block.block_w1_reg\[0\] _03971_ _04315_ sky130_fd_sc_hd__mux2_2
X_15639_ VGND VPWR VGND VPWR _11093_ _11056_ _11097_ _11096_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_29_643 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_115_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_267_1425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_602 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18358_ VPWR VGND VPWR VGND _04253_ block[122] _04213_ enc_block.block_w0_reg\[26\]
+ _04171_ _04254_ sky130_fd_sc_hd__a221o_2
XFILLER_0_28_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_267_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17309_ VGND VPWR VGND VPWR _02701_ _02696_ _03404_ _03403_ sky130_fd_sc_hd__a21oi_2
X_18289_ VPWR VGND VGND VPWR _04191_ _04192_ _04190_ sky130_fd_sc_hd__nor2_2
X_20320_ VGND VPWR VPWR VGND _05580_ _03015_ keymem.key_mem\[9\]\[46\] _05586_ sky130_fd_sc_hd__mux2_2
XFILLER_0_128_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_765 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_124_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_787 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_24_392 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20251_ VGND VPWR VPWR VGND _05546_ _11040_ keymem.key_mem\[9\]\[13\] _05550_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20182_ VGND VPWR _00866_ _05511_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_112_2_Left_583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_177_64 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_50_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24990_ VGND VPWR VPWR VGND clk _01483_ reset_n keymem.key_mem\[5\]\[87\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_239_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23941_ VGND VPWR VPWR VGND clk _00434_ reset_n keymem.key_mem\[13\]\[62\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23872_ VGND VPWR VPWR VGND clk _00365_ reset_n enc_block.block_w2_reg\[25\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_135_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_236_Left_503 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25611_ VGND VPWR VPWR VGND clk _02104_ reset_n keymem.key_mem\[0\]\[68\] sky130_fd_sc_hd__dfrtp_2
X_22823_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[122\] _06839_ _03864_ _05079_ _02158_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_135_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_17_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1070 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_196_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25542_ VGND VPWR VPWR VGND clk _02035_ reset_n keymem.key_mem\[1\]\[127\] sky130_fd_sc_hd__dfrtp_2
X_22754_ VGND VPWR _02107_ _06842_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21705_ VGND VPWR VPWR VGND _06319_ _03099_ keymem.key_mem\[4\]\[55\] _06322_ sky130_fd_sc_hd__mux2_2
X_25473_ VGND VPWR VPWR VGND clk _01966_ reset_n keymem.key_mem\[1\]\[58\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_211_1446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22685_ VGND VPWR _02066_ _06814_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_211_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24424_ VGND VPWR VPWR VGND clk _00917_ reset_n keymem.key_mem\[9\]\[33\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21636_ VGND VPWR _01546_ _06285_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_246_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_62_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24355_ VGND VPWR VPWR VGND clk _00848_ reset_n keymem.key_mem\[10\]\[92\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21567_ VGND VPWR VPWR VGND _06242_ _03613_ keymem.key_mem\[5\]\[119\] _06248_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_245_Left_512 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23306_ VPWR VGND VPWR VGND _07187_ _07185_ _07186_ sky130_fd_sc_hd__or2_2
X_20518_ VGND VPWR VGND VPWR _05676_ _10913_ _01023_ _05690_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_34_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21498_ VGND VPWR VPWR VGND _06209_ _03383_ keymem.key_mem\[5\]\[86\] _06212_ sky130_fd_sc_hd__mux2_2
X_24286_ VGND VPWR VPWR VGND clk _00779_ reset_n keymem.key_mem\[10\]\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_142_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23237_ VPWR VGND _07125_ _07124_ enc_block.round_key\[3\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_20449_ VGND VPWR _00991_ _05653_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_28_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23168_ VGND VPWR VPWR VGND _07054_ _03606_ keymem.prev_key1_reg\[118\] _07069_ sky130_fd_sc_hd__mux2_2
XFILLER_0_100_261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22119_ VGND VPWR VPWR VGND _06538_ _05075_ keymem.key_mem\[3\]\[120\] _06543_ sky130_fd_sc_hd__mux2_2
X_23099_ VGND VPWR VGND VPWR _03431_ _06928_ _03433_ _07026_ sky130_fd_sc_hd__a21o_2
X_15990_ VGND VPWR VGND VPWR _11445_ key[144] _11446_ _11151_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_234_405 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_140_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14941_ VGND VPWR VGND VPWR _10405_ enc_block.sword_ctr_reg\[0\] enc_block.block_w1_reg\[11\]
+ enc_block.sword_ctr_reg\[1\] sky130_fd_sc_hd__and3b_2
XPHY_EDGE_ROW_254_Left_521 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17660_ VGND VPWR _03703_ _03674_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14872_ VPWR VGND VGND VPWR _09122_ _10337_ _09138_ sky130_fd_sc_hd__nor2_2
XFILLER_0_255_1362 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_471 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16611_ VGND VPWR VGND VPWR keymem.rcon_logic.tmp_rcon\[5\] _02458_ _02430_ _02767_
+ sky130_fd_sc_hd__nand3b_2
X_13823_ VPWR VGND VGND VPWR _09294_ _09295_ _09268_ sky130_fd_sc_hd__nor2_2
X_25809_ keymem.prev_key1_reg\[125\] clk _02302_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_138_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17591_ VGND VPWR VGND VPWR _03650_ _02928_ _02877_ key[125] sky130_fd_sc_hd__o21a_2
XFILLER_0_106_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_35_1121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19330_ VGND VPWR _00478_ _05047_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16542_ VPWR VGND VGND VPWR _02700_ _02699_ _07387_ _02697_ _02698_ _02701_ sky130_fd_sc_hd__a311o_2
X_13754_ VGND VPWR VGND VPWR _09080_ _09138_ _09097_ _09127_ _09226_ sky130_fd_sc_hd__a31o_2
XFILLER_0_15_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_188_2_Left_659 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19261_ VGND VPWR _00453_ _05003_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12705_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[54\] _07702_ keymem.key_mem\[2\]\[54\]
+ _07646_ _08254_ sky130_fd_sc_hd__a22o_2
XFILLER_0_6_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16473_ VGND VPWR VGND VPWR _11325_ _11326_ _11275_ _11344_ _02634_ sky130_fd_sc_hd__o22a_2
X_13685_ VGND VPWR _09157_ _09016_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_440 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18212_ VPWR VGND VPWR VGND _04121_ _04045_ _04119_ sky130_fd_sc_hd__or2_2
XFILLER_0_122_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15424_ VPWR VGND VGND VPWR _10475_ _10885_ _10480_ sky130_fd_sc_hd__nor2_2
XFILLER_0_26_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12636_ VGND VPWR enc_block.round_key\[47\] _08191_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19192_ VPWR VGND keymem.key_mem\[13\]\[54\] _04962_ _04961_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_249_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_182_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_65_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18143_ VPWR VGND VPWR VGND _04058_ enc_block.block_w3_reg\[6\] _04056_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_263_Left_530 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15355_ VGND VPWR VPWR VGND _10815_ _10816_ keymem.prev_key0_reg\[106\] _10817_ sky130_fd_sc_hd__or3_2
X_12567_ VGND VPWR VGND VPWR _07877_ keymem.key_mem\[10\]\[41\] _08126_ _08128_ _08129_
+ _08020_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_142_117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_26_679 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_80_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14306_ VPWR VGND VGND VPWR _09476_ _09776_ _09431_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18074_ VPWR VGND VGND VPWR _03994_ _03995_ _03993_ sky130_fd_sc_hd__nor2_2
X_15286_ VGND VPWR _00021_ _10748_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12498_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[35\] _07845_ keymem.key_mem\[2\]\[35\]
+ _07647_ _08066_ sky130_fd_sc_hd__a22o_2
X_17025_ VGND VPWR VGND VPWR _03149_ _11151_ key[188] _03144_ _03148_ sky130_fd_sc_hd__a211o_2
X_14237_ VPWR VGND VGND VPWR _09075_ _09686_ _09697_ _09707_ _09708_ sky130_fd_sc_hd__and4b_2
XFILLER_0_46_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_362 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_238_722 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14168_ VGND VPWR VGND VPWR _09629_ _09589_ keymem.round_ctr_reg\[0\] _09639_ sky130_fd_sc_hd__a21o_2
X_13119_ VGND VPWR VGND VPWR _07648_ keymem.key_mem\[2\]\[95\] _08624_ _08626_ _08627_
+ _08599_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_193_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18976_ VGND VPWR _04809_ enc_block.block_w3_reg\[22\] enc_block.block_w2_reg\[31\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_14099_ VPWR VGND VPWR VGND _09567_ _09569_ _09568_ _09561_ _09570_ sky130_fd_sc_hd__or4_2
XFILLER_0_225_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17927_ VGND VPWR _00240_ _03882_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_56_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17858_ VGND VPWR _03308_ _11044_ _03835_ _03789_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_117_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16809_ VPWR VGND VGND VPWR keylen _02952_ keymem.prev_key1_reg\[40\] _10287_ _10377_
+ _02953_ sky130_fd_sc_hd__a311o_2
XFILLER_0_221_644 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17789_ VGND VPWR VGND VPWR _03736_ keymem.prev_key0_reg\[56\] _03787_ _00197_ sky130_fd_sc_hd__a21o_2
XFILLER_0_117_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19528_ VPWR VGND keymem.key_mem\[12\]\[59\] _05165_ _05158_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_14_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19459_ VGND VPWR VGND VPWR _05127_ keymem.key_mem_we _02765_ _05121_ _00527_ sky130_fd_sc_hd__a31o_2
XFILLER_0_158_283 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_158_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22470_ VGND VPWR _01936_ _06729_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_9_879 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_130_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_133_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21421_ VGND VPWR _01445_ _06171_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_98_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_71_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21352_ VGND VPWR _01412_ _06135_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24140_ VGND VPWR VPWR VGND clk _00633_ reset_n keymem.key_mem\[11\]\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_551 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_128_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20303_ VGND VPWR VPWR VGND _05569_ _02934_ keymem.key_mem\[9\]\[38\] _05577_ sky130_fd_sc_hd__mux2_2
XFILLER_0_13_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_188_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_584 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24071_ VGND VPWR VPWR VGND clk _00564_ reset_n keymem.key_mem\[12\]\[64\] sky130_fd_sc_hd__dfrtp_2
X_21283_ VGND VPWR _01381_ _06097_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_12_340 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_25_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_660 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_141_194 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_229_722 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20234_ VGND VPWR VPWR VGND _05535_ _10194_ keymem.key_mem\[9\]\[5\] _05541_ sky130_fd_sc_hd__mux2_2
XFILLER_0_188_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23022_ VGND VPWR VPWR VGND _02237_ _03144_ _03148_ _06925_ _06980_ sky130_fd_sc_hd__o31a_2
XFILLER_0_25_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1250 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_198_1338 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_99_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20165_ VGND VPWR _00858_ _05502_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_31_Left_299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_99_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20096_ VGND VPWR _00825_ _05466_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24973_ VGND VPWR VPWR VGND clk _01466_ reset_n keymem.key_mem\[5\]\[70\] sky130_fd_sc_hd__dfrtp_2
X_23924_ VGND VPWR VPWR VGND clk _00417_ reset_n keymem.key_mem\[13\]\[45\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_97_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23855_ VGND VPWR VPWR VGND clk _00348_ reset_n enc_block.block_w2_reg\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_1176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_139_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_170_1235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22806_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[107\] _06858_ _06857_ _05048_ _02143_
+ sky130_fd_sc_hd__a22o_2
X_23786_ VGND VPWR VPWR VGND clk _00279_ reset_n enc_block.block_w0_reg\[5\] sky130_fd_sc_hd__dfrtp_2
X_20998_ VGND VPWR VPWR VGND _05945_ _05048_ keymem.key_mem\[7\]\[107\] _05947_ sky130_fd_sc_hd__mux2_2
XFILLER_0_36_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25525_ VGND VPWR VPWR VGND clk _02018_ reset_n keymem.key_mem\[1\]\[110\] sky130_fd_sc_hd__dfrtp_2
X_22737_ VGND VPWR VPWR VGND _06833_ keymem.key_mem\[0\]\[63\] _03184_ _06834_ sky130_fd_sc_hd__mux2_2
XFILLER_0_109_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_48_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13470_ VGND VPWR _08942_ _08941_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25456_ VGND VPWR VPWR VGND clk _01949_ reset_n keymem.key_mem\[1\]\[41\] sky130_fd_sc_hd__dfrtp_2
X_22668_ VGND VPWR _02058_ _06805_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_211_1298 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_47_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_246_1317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12421_ VPWR VGND VPWR VGND _07995_ keymem.key_mem\[5\]\[28\] _07613_ keymem.key_mem\[8\]\[28\]
+ _07903_ _07996_ sky130_fd_sc_hd__a221o_2
X_24407_ VGND VPWR VPWR VGND clk _00900_ reset_n keymem.key_mem\[9\]\[16\] sky130_fd_sc_hd__dfrtp_2
X_21619_ VGND VPWR VPWR VGND _06275_ _11098_ keymem.key_mem\[4\]\[14\] _06277_ sky130_fd_sc_hd__mux2_2
X_25387_ VGND VPWR VPWR VGND clk _01880_ reset_n keymem.key_mem\[2\]\[100\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_168_1164 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_465 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_62_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22599_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[111\] _06775_ _06774_ _05056_ _02019_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_1_1472 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15140_ VGND VPWR _10604_ _10603_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_63_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24338_ VGND VPWR VPWR VGND clk _00831_ reset_n keymem.key_mem\[10\]\[75\] sky130_fd_sc_hd__dfrtp_2
X_12352_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[21\] _07535_ _07933_ _07928_ _07934_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_181_1320 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_284 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_146_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15071_ VGND VPWR _10535_ _10534_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_50_457 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_65_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_107_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12283_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[16\] _07535_ _07869_ _07864_ _07870_
+ sky130_fd_sc_hd__o22a_2
X_24269_ VGND VPWR VPWR VGND clk _00762_ reset_n keymem.key_mem\[10\]\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_43_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14022_ VGND VPWR VPWR VGND _09304_ _09317_ _09303_ _09494_ sky130_fd_sc_hd__or3_2
XFILLER_0_107_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_356 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18830_ _04676_ _04678_ _03982_ _04677_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_248_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_257_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18761_ VPWR VGND _04615_ enc_block.block_w2_reg\[26\] enc_block.block_w3_reg\[18\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_15973_ _11340_ _11429_ _11391_ _11408_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_257_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14924_ enc_block.sword_ctr_reg\[1\] _10388_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[9\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_17712_ VGND VPWR VGND VPWR _03732_ keymem.prev_key1_reg\[26\] _03741_ _03733_ sky130_fd_sc_hd__a21oi_2
X_18692_ VGND VPWR _04553_ _04496_ _04552_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_250_728 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_264_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17643_ VGND VPWR _03691_ _03211_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_118_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14855_ VGND VPWR VPWR VGND _09927_ _10319_ key[135] _10320_ sky130_fd_sc_hd__mux2_2
X_13806_ VGND VPWR VGND VPWR enc_block.block_w1_reg\[30\] _08948_ _09022_ _09276_
+ _09278_ _09277_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_118_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_54_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17574_ VPWR VGND VGND VPWR _03635_ _03240_ _02750_ sky130_fd_sc_hd__nand2_2
X_14786_ VGND VPWR VGND VPWR _09293_ _09403_ _09323_ _09449_ _10252_ sky130_fd_sc_hd__o22a_2
X_11998_ VPWR VGND VGND VPWR _07532_ _07601_ _07530_ sky130_fd_sc_hd__nor2_2
XFILLER_0_15_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19313_ VGND VPWR VPWR VGND _05025_ _05035_ keymem.key_mem\[13\]\[101\] _05036_ sky130_fd_sc_hd__mux2_2
XFILLER_0_188_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16525_ VGND VPWR VGND VPWR _02682_ _02681_ _02685_ _02683_ sky130_fd_sc_hd__a21oi_2
X_13737_ VGND VPWR VGND VPWR _09209_ _09065_ _09051_ _09057_ _09010_ sky130_fd_sc_hd__a211o_2
XFILLER_0_133_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16456_ VPWR VGND VPWR VGND _02452_ _02348_ _02617_ _11579_ _02438_ sky130_fd_sc_hd__or4b_2
X_19244_ VPWR VGND keymem.key_mem_we _04992_ _03295_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_27_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13668_ VGND VPWR _09140_ _09139_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_160_2_Right_232 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_186_1220 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15407_ VPWR VGND VGND VPWR _10867_ _10530_ _10546_ _10543_ _10868_ _10580_ sky130_fd_sc_hd__o221a_2
X_12619_ VPWR VGND VPWR VGND _08175_ keymem.key_mem\[13\]\[46\] _07731_ keymem.key_mem\[14\]\[46\]
+ _07721_ _08176_ sky130_fd_sc_hd__a221o_2
XFILLER_0_229_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19175_ VGND VPWR _04951_ _04876_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_186_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16387_ VGND VPWR _02550_ _02549_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13599_ VPWR VGND VGND VPWR _09071_ _09057_ _09058_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18126_ VPWR VGND VGND VPWR _04042_ _04043_ _04041_ sky130_fd_sc_hd__nor2_2
XFILLER_0_108_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15338_ VGND VPWR VGND VPWR _10547_ _10667_ _10574_ _10800_ sky130_fd_sc_hd__a21o_2
XFILLER_0_206_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_638 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_252_Right_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_130_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_278 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18057_ VGND VPWR _03978_ _03977_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15269_ VGND VPWR _10732_ _09987_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_123_172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_125_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_183 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17008_ VGND VPWR VPWR VGND _11109_ _03132_ key[59] _03133_ sky130_fd_sc_hd__mux2_2
XFILLER_0_50_991 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_205_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_111_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_201_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_899 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18959_ VPWR VGND VGND VPWR _04793_ _04794_ _04382_ sky130_fd_sc_hd__nor2_2
XFILLER_0_253_555 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21970_ VGND VPWR _01701_ _06464_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_20_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_471 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_154_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20921_ VGND VPWR _01210_ _05906_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_90_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_94_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_441 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23640_ VPWR VGND VPWR VGND keymem.key_mem_ctrl_reg\[0\] reset_n _00009_ clk sky130_fd_sc_hd__dfstp_2
X_20852_ VGND VPWR VPWR VGND _05867_ _04931_ keymem.key_mem\[7\]\[38\] _05870_ sky130_fd_sc_hd__mux2_2
XFILLER_0_7_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23571_ VGND VPWR VPWR VGND clk _00072_ reset_n keymem.key_mem\[14\]\[60\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_212_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20783_ VGND VPWR VGND VPWR _05832_ keymem.key_mem_we _10284_ _05821_ _01146_ sky130_fd_sc_hd__a31o_2
XFILLER_0_64_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25310_ VGND VPWR VPWR VGND clk _01803_ reset_n keymem.key_mem\[2\]\[23\] sky130_fd_sc_hd__dfrtp_2
X_22522_ VGND VPWR _01969_ _06748_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_130_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1030 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25241_ VGND VPWR VPWR VGND clk _01734_ reset_n keymem.key_mem\[3\]\[82\] sky130_fd_sc_hd__dfrtp_2
X_22453_ VGND VPWR _01928_ _06720_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_267_1074 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_31_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_146_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_267_1096 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21404_ VGND VPWR VPWR VGND _06162_ _02964_ keymem.key_mem\[5\]\[41\] _06163_ sky130_fd_sc_hd__mux2_2
XFILLER_0_44_273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25172_ VGND VPWR VPWR VGND clk _01665_ reset_n keymem.key_mem\[3\]\[13\] sky130_fd_sc_hd__dfrtp_2
X_22384_ VGND VPWR _01896_ _06683_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_165_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24123_ VGND VPWR VPWR VGND clk _00616_ reset_n keymem.key_mem\[12\]\[116\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_370 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21335_ VGND VPWR _01404_ _06126_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_20_619 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_980 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24054_ VGND VPWR VPWR VGND clk _00547_ reset_n keymem.key_mem\[12\]\[47\] sky130_fd_sc_hd__dfrtp_2
X_21266_ VGND VPWR VPWR VGND _06087_ _03525_ keymem.key_mem\[6\]\[105\] _06089_ sky130_fd_sc_hd__mux2_2
XFILLER_0_198_1124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23005_ VGND VPWR _02230_ _06970_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20217_ VGND VPWR _00883_ _05529_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21197_ VGND VPWR VPWR VGND _06052_ _03259_ keymem.key_mem\[6\]\[72\] _06053_ sky130_fd_sc_hd__mux2_2
XFILLER_0_229_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20148_ VGND VPWR VPWR VGND _05493_ _03452_ keymem.key_mem\[10\]\[94\] _05494_ sky130_fd_sc_hd__mux2_2
XFILLER_0_239_1121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_107_1_Left_374 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_102_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20079_ VGND VPWR VPWR VGND _05457_ _03162_ keymem.key_mem\[10\]\[61\] _05458_ sky130_fd_sc_hd__mux2_2
X_24956_ VGND VPWR VPWR VGND clk _01449_ reset_n keymem.key_mem\[5\]\[53\] sky130_fd_sc_hd__dfrtp_2
X_12970_ VPWR VGND VPWR VGND _08492_ keymem.key_mem\[8\]\[80\] _07752_ keymem.key_mem\[1\]\[80\]
+ _07799_ _08493_ sky130_fd_sc_hd__a221o_2
X_11921_ VGND VPWR result[127] _07524_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23907_ VGND VPWR VPWR VGND clk _00400_ reset_n keymem.key_mem\[13\]\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_176_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_213_953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24887_ VGND VPWR VPWR VGND clk _01380_ reset_n keymem.key_mem\[6\]\[112\] sky130_fd_sc_hd__dfrtp_2
X_14640_ VPWR VGND VPWR VGND _10106_ _10107_ _10061_ _10104_ sky130_fd_sc_hd__or3b_2
X_11852_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[29\] dec_new_block\[93\]
+ _07490_ sky130_fd_sc_hd__mux2_2
X_23838_ VGND VPWR VPWR VGND clk _00331_ reset_n enc_block.block_w1_reg\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_213_1338 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_79_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14571_ VGND VPWR VGND VPWR _10038_ _10037_ _10039_ _10036_ _10035_ sky130_fd_sc_hd__nand4_2
X_11783_ VGND VPWR result[58] _07455_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23769_ keymem.prev_key0_reg\[125\] clk _00266_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_55_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_196_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16310_ VGND VPWR VGND VPWR _09511_ _02472_ _02470_ _02471_ _02474_ sky130_fd_sc_hd__a31o_2
X_13522_ VPWR VGND VPWR VGND _08993_ _08985_ _08992_ _08945_ enc_block.block_w2_reg\[4\]
+ _08994_ sky130_fd_sc_hd__a221o_2
X_25508_ VGND VPWR VPWR VGND clk _02001_ reset_n keymem.key_mem\[1\]\[93\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_184_359 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17290_ VPWR VGND VGND VPWR _03386_ _03387_ keylen sky130_fd_sc_hd__nor2_2
XFILLER_0_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_324 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16241_ VGND VPWR VGND VPWR _02405_ key[147] _02406_ _09868_ sky130_fd_sc_hd__a21bo_2
X_25439_ VGND VPWR VPWR VGND clk _01932_ reset_n keymem.key_mem\[1\]\[24\] sky130_fd_sc_hd__dfrtp_2
X_13453_ VGND VPWR _08925_ _08924_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_196_Left_463 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12404_ VPWR VGND VPWR VGND _07980_ keymem.key_mem\[5\]\[26\] _07596_ keymem.key_mem\[13\]\[26\]
+ _07587_ _07981_ sky130_fd_sc_hd__a221o_2
XFILLER_0_35_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16172_ VPWR VGND VGND VPWR _02338_ _02337_ _11623_ _09931_ _09930_ key[18] sky130_fd_sc_hd__o2111a_2
XFILLER_0_10_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13384_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[121\] _08027_ _08865_ _08861_ _08866_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_183_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15123_ VGND VPWR _10587_ _10586_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12335_ VGND VPWR _07918_ _07591_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_50_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15054_ VPWR VGND VPWR VGND _10483_ _10466_ _10453_ _10451_ _10518_ sky130_fd_sc_hd__or4_2
X_19931_ VGND VPWR VPWR VGND _05372_ keymem.key_mem\[11\]\[121\] _03627_ _05378_ sky130_fd_sc_hd__mux2_2
X_12266_ VGND VPWR _07854_ _07551_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_142_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14005_ VPWR VGND VGND VPWR _09401_ _09475_ _09477_ _09410_ _09476_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_142_1178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19862_ VGND VPWR VPWR VGND _05339_ keymem.key_mem\[11\]\[88\] _03401_ _05342_ sky130_fd_sc_hd__mux2_2
XFILLER_0_120_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12197_ VPWR VGND VPWR VGND keymem.key_mem\[4\]\[10\] _07692_ keymem.key_mem\[1\]\[10\]
+ _07714_ _07790_ sky130_fd_sc_hd__a22o_2
X_18813_ VPWR VGND _04663_ _04662_ enc_block.round_key\[38\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_120_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19793_ VGND VPWR VPWR VGND _05303_ keymem.key_mem\[11\]\[55\] _03099_ _05306_ sky130_fd_sc_hd__mux2_2
XFILLER_0_120_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18744_ VGND VPWR _04600_ _04599_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_235_577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_194_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15956_ VPWR VGND VGND VPWR _11221_ _11412_ _11286_ sky130_fd_sc_hd__nor2_2
XFILLER_0_204_920 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_190_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14907_ VGND VPWR _10371_ _09732_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15887_ VPWR VGND VPWR VGND _11206_ _11202_ _11207_ _11187_ _11343_ sky130_fd_sc_hd__or4_2
X_18675_ VGND VPWR _04538_ _04536_ _04537_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_91_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_144_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17626_ VGND VPWR _03679_ _03211_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_156_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14838_ VPWR VGND VPWR VGND _09448_ _10302_ _10301_ _10300_ _10303_ sky130_fd_sc_hd__or4_2
XFILLER_0_187_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1079 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_59_866 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14769_ VPWR VGND VPWR VGND _09567_ _09735_ _09584_ _10234_ _10235_ sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_69_2_Left_540 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17557_ VGND VPWR VPWR VGND _03593_ keymem.key_mem\[14\]\[120\] _03620_ _03621_ sky130_fd_sc_hd__mux2_2
XFILLER_0_59_888 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_187_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_175_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_58_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16508_ VGND VPWR VGND VPWR _11438_ _11301_ _02668_ keymem.rcon_reg\[0\] sky130_fd_sc_hd__a21oi_2
XFILLER_0_89_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17488_ VGND VPWR VPWR VGND _03534_ keymem.key_mem\[14\]\[111\] _03560_ _03561_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_121_2_Left_592 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_128_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_131_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_190_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19227_ VPWR VGND keymem.key_mem\[13\]\[69\] _04982_ _04979_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16439_ VPWR VGND VPWR VGND keymem.prev_key1_reg\[54\] _02601_ _02599_ _02600_ sky130_fd_sc_hd__or3b_2
XPHY_EDGE_ROW_161_2_Right_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_61_519 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_27_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19158_ VGND VPWR VPWR VGND _04928_ _04939_ keymem.key_mem\[13\]\[42\] _04940_ sky130_fd_sc_hd__mux2_2
X_18109_ VPWR VGND VGND VPWR _04026_ _04027_ _03966_ sky130_fd_sc_hd__nor2_2
X_19089_ VPWR VGND keymem.key_mem\[13\]\[14\] _04899_ _04887_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_2_852 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_200_Left_467 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_257_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21120_ VGND VPWR _01303_ _06012_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_172_1_Left_439 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_78_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_246_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_199_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_850 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_239_861 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21051_ VGND VPWR VPWR VGND _05972_ _09991_ keymem.key_mem\[6\]\[3\] _05976_ sky130_fd_sc_hd__mux2_2
XFILLER_0_240_1291 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20002_ VGND VPWR _00780_ _05417_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_254_831 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_185_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_201_1275 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24810_ VGND VPWR VPWR VGND clk _01303_ reset_n keymem.key_mem\[6\]\[35\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25790_ keymem.prev_key1_reg\[106\] clk _02283_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_24741_ VGND VPWR VPWR VGND clk _01234_ reset_n keymem.key_mem\[7\]\[94\] sky130_fd_sc_hd__dfrtp_2
X_21953_ VGND VPWR _01693_ _06455_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_234_1040 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_178_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_55_1146 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_94_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20904_ VGND VPWR VGND VPWR _05897_ keymem.key_mem_we _03173_ _05893_ _01202_ sky130_fd_sc_hd__a31o_2
X_24672_ VGND VPWR VPWR VGND clk _01165_ reset_n keymem.key_mem\[7\]\[25\] sky130_fd_sc_hd__dfrtp_2
X_21884_ VPWR VGND keymem.key_mem\[3\]\[10\] _06418_ _06413_ VPWR VGND sky130_fd_sc_hd__and2_2
X_23623_ VGND VPWR VPWR VGND clk _00124_ reset_n keymem.key_mem\[14\]\[112\] sky130_fd_sc_hd__dfrtp_2
X_20835_ VGND VPWR VGND VPWR _05860_ keymem.key_mem_we _02839_ _05850_ _01170_ sky130_fd_sc_hd__a31o_2
XFILLER_0_204_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23554_ VGND VPWR VPWR VGND clk _00055_ reset_n keymem.key_mem\[14\]\[43\] sky130_fd_sc_hd__dfrtp_2
X_20766_ VPWR VGND VPWR VGND _05822_ keymem.round_ctr_reg\[3\] _05818_ sky130_fd_sc_hd__or2_2
XFILLER_0_247_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22505_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[52\] _06737_ _06736_ _04958_ _01960_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_52_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23485_ VPWR VGND VPWR VGND _07346_ block[29] _03958_ enc_block.block_w3_reg\[29\]
+ _04504_ _07347_ sky130_fd_sc_hd__a221o_2
X_20697_ VGND VPWR _01108_ _05784_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_18_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25224_ VGND VPWR VPWR VGND clk _01717_ reset_n keymem.key_mem\[3\]\[65\] sky130_fd_sc_hd__dfrtp_2
X_22436_ VGND VPWR _01920_ _06711_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_208_1418 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_208_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_134_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25155_ VGND VPWR VPWR VGND clk _01648_ reset_n keymem.key_mem\[4\]\[124\] sky130_fd_sc_hd__dfrtp_2
X_22367_ VGND VPWR _01888_ _06674_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_32_265 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12120_ VGND VPWR _07717_ _07716_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24106_ VGND VPWR VPWR VGND clk _00599_ reset_n keymem.key_mem\[12\]\[99\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_108_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21318_ VGND VPWR VPWR VGND _06117_ _09536_ keymem.key_mem\[5\]\[0\] _06118_ sky130_fd_sc_hd__mux2_2
X_25086_ VGND VPWR VPWR VGND clk _01579_ reset_n keymem.key_mem\[4\]\[55\] sky130_fd_sc_hd__dfrtp_2
X_22298_ VGND VPWR _06638_ _03287_ _01855_ _06567_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_206_1175 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12051_ VGND VPWR _07651_ _07602_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24037_ VGND VPWR VPWR VGND clk _00530_ reset_n keymem.key_mem\[12\]\[30\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_186 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21249_ VGND VPWR VPWR VGND _06076_ _03474_ keymem.key_mem\[6\]\[97\] _06080_ sky130_fd_sc_hd__mux2_2
XFILLER_0_263_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_229_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_229_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_258_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_555 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15810_ VGND VPWR _11266_ _11265_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_219_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16790_ VGND VPWR _00050_ _02935_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_245_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15741_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[20\] _10402_ _11197_ _09255_ _11195_
+ _11196_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_219_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12953_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[79\] _07652_ keymem.key_mem\[11\]\[79\]
+ _07809_ _08477_ sky130_fd_sc_hd__a22o_2
X_24939_ VGND VPWR VPWR VGND clk _01432_ reset_n keymem.key_mem\[5\]\[36\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_137_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11904_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[23\] dec_new_block\[119\]
+ _07516_ sky130_fd_sc_hd__mux2_2
XFILLER_0_73_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_440 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15672_ VGND VPWR VPWR VGND _10751_ _10668_ _11129_ _11128_ _11127_ sky130_fd_sc_hd__o211a_2
X_18460_ VPWR VGND VPWR VGND _04345_ _04341_ _04344_ sky130_fd_sc_hd__or2_2
X_12884_ VPWR VGND VPWR VGND _08414_ keymem.key_mem\[14\]\[72\] _07666_ keymem.key_mem\[10\]\[72\]
+ _07876_ _08415_ sky130_fd_sc_hd__a221o_2
XFILLER_0_154_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_73_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17411_ VGND VPWR _03494_ _02866_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_157_315 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14623_ VGND VPWR _10091_ _09511_ VPWR VGND sky130_fd_sc_hd__buf_1
X_11835_ VGND VPWR result[84] _07481_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18391_ VPWR VGND VGND VPWR _04283_ _04284_ _04190_ sky130_fd_sc_hd__nor2_2
XFILLER_0_200_455 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_67_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17342_ VPWR VGND VPWR VGND _03433_ _02677_ _03431_ key[220] _10838_ _03434_ sky130_fd_sc_hd__a221o_2
X_14554_ VPWR VGND VPWR VGND _10022_ _09937_ _10021_ sky130_fd_sc_hd__or2_2
XFILLER_0_200_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11766_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[18\] dec_new_block\[50\]
+ _07447_ sky130_fd_sc_hd__mux2_2
XFILLER_0_56_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13505_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[7\] _08956_ _08977_ _08943_ _08975_
+ _08976_ sky130_fd_sc_hd__a32oi_2
X_17273_ VPWR VGND VGND VPWR _03372_ key[213] _03077_ sky130_fd_sc_hd__nand2_2
XFILLER_0_113_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14485_ VPWR VGND VPWR VGND _09949_ _09953_ _09951_ _09947_ _09954_ sky130_fd_sc_hd__or4_2
XFILLER_0_99_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11697_ VGND VPWR result[15] _07412_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16224_ VGND VPWR VGND VPWR _11239_ _11466_ _11284_ _11367_ _02389_ sky130_fd_sc_hd__o22a_2
XFILLER_0_10_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19012_ VPWR VGND VPWR VGND _04841_ _04625_ _04839_ sky130_fd_sc_hd__or2_2
X_13436_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[127\] _07652_ keymem.key_mem\[4\]\[127\]
+ _07914_ _08912_ sky130_fd_sc_hd__a22o_2
XFILLER_0_183_1223 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_183_1234 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_51_530 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_84_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16155_ VGND VPWR VGND VPWR _11609_ _11417_ _11291_ _11230_ _11564_ _11412_ sky130_fd_sc_hd__a32o_2
XFILLER_0_148_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13367_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[120\] _07742_ keymem.key_mem\[12\]\[120\]
+ _07620_ _08850_ sky130_fd_sc_hd__a22o_2
XFILLER_0_267_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15106_ VPWR VGND VGND VPWR _10485_ _10569_ _10570_ _10513_ _10519_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_45_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12318_ VGND VPWR _07902_ _07861_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_80_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16086_ VGND VPWR VGND VPWR _11539_ _11538_ _11541_ _11540_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_267_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13298_ VPWR VGND VPWR VGND _08787_ keymem.key_mem\[12\]\[113\] _07807_ keymem.key_mem\[8\]\[113\]
+ _07929_ _08788_ sky130_fd_sc_hd__a221o_2
XFILLER_0_20_950 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15037_ VGND VPWR VGND VPWR _10501_ _10500_ _10472_ _10440_ _10464_ sky130_fd_sc_hd__a211o_2
XFILLER_0_255_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19914_ VGND VPWR VPWR VGND _05361_ keymem.key_mem\[11\]\[113\] _03573_ _05369_ sky130_fd_sc_hd__mux2_2
X_12249_ VGND VPWR _07838_ _07761_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_267_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_500 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1083 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19845_ VGND VPWR VPWR VGND _05328_ keymem.key_mem\[11\]\[80\] _03330_ _05333_ sky130_fd_sc_hd__mux2_2
XFILLER_0_120_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19776_ VGND VPWR VPWR VGND _05292_ keymem.key_mem\[11\]\[47\] _03025_ _05297_ sky130_fd_sc_hd__mux2_2
XFILLER_0_21_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_834 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16988_ VGND VPWR VGND VPWR _02713_ _02712_ _03115_ keymem.prev_key1_reg\[57\] sky130_fd_sc_hd__a21oi_2
XFILLER_0_257_1073 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18727_ VGND VPWR _04584_ enc_block.block_w0_reg\[7\] _04383_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_251_856 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_262_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15939_ VGND VPWR _11395_ _11180_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_95_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_155_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_889 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18658_ VPWR VGND VPWR VGND _04523_ _04307_ _04522_ sky130_fd_sc_hd__or2_2
XFILLER_0_56_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_203_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17609_ VPWR VGND VGND VPWR _11456_ _03666_ key[255] sky130_fd_sc_hd__nor2_2
X_18589_ VPWR VGND _04461_ enc_block.block_w0_reg\[0\] enc_block.block_w2_reg\[23\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_4_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20620_ VGND VPWR VPWR VGND _05736_ _03149_ keymem.key_mem\[8\]\[60\] _05744_ sky130_fd_sc_hd__mux2_2
XFILLER_0_19_538 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_188_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_188_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_944 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_131_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20551_ VGND VPWR VPWR VGND _05703_ _02764_ keymem.key_mem\[8\]\[27\] _05708_ sky130_fd_sc_hd__mux2_2
XFILLER_0_6_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23270_ VPWR VGND _07155_ _07154_ enc_block.round_key\[6\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_89_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_162_2_Right_234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20482_ VGND VPWR _01007_ _05670_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_116_278 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_80_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_162_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22221_ VGND VPWR VPWR VGND _06589_ _02945_ keymem.key_mem\[2\]\[39\] _06598_ sky130_fd_sc_hd__mux2_2
XFILLER_0_166_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22152_ VGND VPWR _01786_ _06561_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21103_ VGND VPWR _01295_ _06003_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_196_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_258_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22083_ VGND VPWR VPWR VGND _06516_ _05039_ keymem.key_mem\[3\]\[103\] _06524_ sky130_fd_sc_hd__mux2_2
XFILLER_0_61_1172 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21034_ VGND VPWR _01264_ _05965_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_103_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_201_1061 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_129_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25842_ VGND VPWR VPWR VGND clk _02335_ reset_n enc_block.block_w3_reg\[30\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_236_1102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25773_ keymem.prev_key1_reg\[89\] clk _02266_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22985_ VGND VPWR VGND VPWR _02222_ _06958_ _06954_ keymem.prev_key1_reg\[45\] sky130_fd_sc_hd__o21a_2
XFILLER_0_173_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24724_ VGND VPWR VPWR VGND clk _01217_ reset_n keymem.key_mem\[7\]\[77\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_74_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21936_ VGND VPWR _06446_ _06403_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_214_1422 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24655_ VGND VPWR VPWR VGND clk _01148_ reset_n keymem.key_mem\[7\]\[8\] sky130_fd_sc_hd__dfrtp_2
X_21867_ VPWR VGND keymem.key_mem\[3\]\[2\] _06409_ _06406_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_139_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23606_ VGND VPWR VPWR VGND clk _00107_ reset_n keymem.key_mem\[14\]\[95\] sky130_fd_sc_hd__dfrtp_2
X_20818_ VGND VPWR VGND VPWR _05851_ keymem.key_mem_we _02608_ _05850_ _01162_ sky130_fd_sc_hd__a31o_2
X_24586_ VGND VPWR VPWR VGND clk _01079_ reset_n keymem.key_mem\[8\]\[67\] sky130_fd_sc_hd__dfrtp_2
X_21798_ VGND VPWR _01623_ _06370_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_38_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_110_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_817 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23537_ VGND VPWR VPWR VGND clk _00038_ reset_n keymem.key_mem\[14\]\[26\] sky130_fd_sc_hd__dfrtp_2
X_20749_ VGND VPWR _01133_ _05811_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_52_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_1537 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_110_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14270_ VPWR VGND VPWR VGND _09740_ _09323_ _09440_ sky130_fd_sc_hd__or2_2
X_23468_ VPWR VGND VPWR VGND _07331_ block[27] _04139_ enc_block.block_w3_reg\[27\]
+ _04138_ _07332_ sky130_fd_sc_hd__a221o_2
XFILLER_0_184_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_530 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25207_ VGND VPWR VPWR VGND clk _01700_ reset_n keymem.key_mem\[3\]\[48\] sky130_fd_sc_hd__dfrtp_2
X_13221_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[105\] _07748_ keymem.key_mem\[1\]\[105\]
+ _07558_ _08719_ sky130_fd_sc_hd__a22o_2
XFILLER_0_180_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_243_1128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_247_1297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22419_ VGND VPWR VPWR VGND _06702_ keymem.key_mem\[1\]\[4\] _10099_ _06703_ sky130_fd_sc_hd__mux2_2
X_23399_ VGND VPWR VGND VPWR _07270_ _04505_ _07268_ _07269_ _07271_ sky130_fd_sc_hd__a31o_2
XFILLER_0_81_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_33_596 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13152_ VPWR VGND VPWR VGND _08656_ keymem.key_mem\[8\]\[98\] _07541_ keymem.key_mem\[4\]\[98\]
+ _07854_ _08657_ sky130_fd_sc_hd__a221o_2
X_25138_ VGND VPWR VPWR VGND clk _01631_ reset_n keymem.key_mem\[4\]\[107\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_260_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1404 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_758 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12103_ VGND VPWR VGND VPWR _07691_ keymem.key_mem\[3\]\[5\] _07696_ _07700_ _07701_
+ _07663_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_130_270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17960_ VGND VPWR VPWR VGND _03896_ _03904_ keymem.prev_key0_reg\[110\] _03905_ sky130_fd_sc_hd__mux2_2
X_13083_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[91\] _08577_ _08594_ _08590_ _08595_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_260_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25069_ VGND VPWR VPWR VGND clk _01562_ reset_n keymem.key_mem\[4\]\[38\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_40_1201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16911_ VPWR VGND VPWR VGND _03045_ _03038_ _03037_ key[177] _03027_ _03046_ sky130_fd_sc_hd__a221o_2
X_12034_ VGND VPWR VGND VPWR _07629_ keymem.key_mem\[10\]\[2\] _07630_ _07634_ _07635_
+ _07616_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_109_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17891_ VGND VPWR VPWR VGND _03729_ _03857_ _03399_ _03858_ sky130_fd_sc_hd__or3_2
XFILLER_0_40_1256 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_121_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_864 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19630_ VGND VPWR _00607_ _05218_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_178_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16842_ VPWR VGND VGND VPWR _02983_ _02978_ _02981_ sky130_fd_sc_hd__nand2_2
XFILLER_0_256_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_191_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19561_ VPWR VGND VGND VPWR _05182_ keymem.key_mem\[12\]\[75\] _05095_ sky130_fd_sc_hd__nand2_2
X_13985_ VPWR VGND VGND VPWR _09456_ _09457_ _09302_ sky130_fd_sc_hd__nor2_2
X_16773_ VGND VPWR _09931_ key[37] _02920_ _10327_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_191_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_889 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18512_ VGND VPWR _04392_ enc_block.block_w2_reg\[16\] enc_block.block_w1_reg\[24\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_1190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15724_ VGND VPWR _11180_ _11179_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12936_ VGND VPWR VGND VPWR _08008_ keymem.key_mem\[2\]\[77\] _08459_ _08461_ _08462_
+ _07896_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_125_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19492_ VGND VPWR _00542_ _05145_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_232_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_157_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18443_ VPWR VGND VPWR VGND _04329_ _04291_ _04327_ enc_block.block_w1_reg\[1\] _04317_
+ _00309_ sky130_fd_sc_hd__a221o_2
X_15655_ VPWR VGND VPWR VGND _10931_ _10988_ _10980_ _10926_ _11112_ sky130_fd_sc_hd__or4_2
X_12867_ VPWR VGND VPWR VGND keymem.key_mem\[8\]\[70\] _07878_ keymem.key_mem\[1\]\[70\]
+ _07969_ _08400_ sky130_fd_sc_hd__a22o_2
XFILLER_0_201_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_292 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_232_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14606_ VGND VPWR VGND VPWR _10074_ _09888_ _09368_ _10072_ _10073_ sky130_fd_sc_hd__a211o_2
X_11818_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[12\] dec_new_block\[76\]
+ _07473_ sky130_fd_sc_hd__mux2_2
X_18374_ VPWR VGND _04268_ _04021_ enc_block.block_w1_reg\[20\] VPWR VGND sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_89_1_Right_690 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15586_ VPWR VGND VPWR VGND _11044_ keymem.prev_key1_reg\[78\] sky130_fd_sc_hd__inv_2
XFILLER_0_201_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12798_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[63\] _07568_ keymem.key_mem\[8\]\[63\]
+ _07540_ _08338_ sky130_fd_sc_hd__a22o_2
X_14537_ VGND VPWR VGND VPWR _10005_ _09149_ _09100_ _09154_ _09107_ _10004_ sky130_fd_sc_hd__o221ai_2
X_17325_ VGND VPWR VPWR VGND _03384_ keymem.key_mem\[14\]\[90\] _03418_ _03419_ sky130_fd_sc_hd__mux2_2
X_11749_ VGND VPWR result[41] _07438_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_43_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1331 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14468_ VPWR VGND VGND VPWR _09168_ _09937_ _09091_ sky130_fd_sc_hd__nor2_2
XFILLER_0_119_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17256_ VGND VPWR VPWR VGND _03296_ keymem.key_mem\[14\]\[83\] _03356_ _03357_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_113_204 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16207_ VGND VPWR VGND VPWR _02355_ _02371_ _02372_ _02350_ _02363_ sky130_fd_sc_hd__nor4_2
X_13419_ VGND VPWR VGND VPWR _07800_ keymem.key_mem\[1\]\[125\] _08894_ _08896_ _08897_
+ _07573_ sky130_fd_sc_hd__a2111o_2
X_17187_ VPWR VGND VPWR VGND _03294_ _03293_ _03291_ _02497_ _03290_ _03295_ sky130_fd_sc_hd__a221o_2
XFILLER_0_10_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1270 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14399_ VGND VPWR _09868_ _09521_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_148_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_52_894 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16138_ VPWR VGND VGND VPWR _11235_ _11370_ _11592_ _11182_ _11404_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_84_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1009 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_11_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16069_ VGND VPWR VGND VPWR _11376_ _11211_ _11400_ _11283_ _11524_ sky130_fd_sc_hd__o22a_2
XFILLER_0_121_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_267_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_791 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_264_981 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19828_ VGND VPWR VPWR VGND _05314_ keymem.key_mem\[11\]\[72\] _03259_ _05324_ sky130_fd_sc_hd__mux2_2
XFILLER_0_196_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_209_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19759_ VGND VPWR VPWR VGND _05281_ keymem.key_mem\[11\]\[39\] _02945_ _05288_ sky130_fd_sc_hd__mux2_2
XFILLER_0_159_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22770_ VGND VPWR _02118_ _06847_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_155_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21721_ VGND VPWR _06330_ _06262_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_8_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24440_ VGND VPWR VPWR VGND clk _00933_ reset_n keymem.key_mem\[9\]\[49\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_231_1065 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21652_ VGND VPWR VPWR VGND _06286_ _02838_ keymem.key_mem\[4\]\[30\] _06294_ sky130_fd_sc_hd__mux2_2
XFILLER_0_93_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20603_ VGND VPWR VPWR VGND _05725_ _03075_ keymem.key_mem\[8\]\[52\] _05735_ sky130_fd_sc_hd__mux2_2
XFILLER_0_35_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24371_ VGND VPWR VPWR VGND clk _00864_ reset_n keymem.key_mem\[10\]\[108\] sky130_fd_sc_hd__dfrtp_2
X_21583_ VGND VPWR VPWR VGND _06116_ _03668_ keymem.key_mem\[5\]\[127\] _06256_ sky130_fd_sc_hd__mux2_2
XFILLER_0_163_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23322_ VGND VPWR VGND VPWR _07201_ _04266_ _07095_ _07202_ enc_block.block_w3_reg\[11\]
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_34_338 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_209_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20534_ VGND VPWR VPWR VGND _05692_ _02409_ keymem.key_mem\[8\]\[19\] _05699_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_116_1_Left_383 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_7_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_166_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23253_ VGND VPWR _02309_ _07139_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_163_2_Right_235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_127_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20465_ VGND VPWR VPWR VGND _05660_ _03585_ keymem.key_mem\[9\]\[115\] _05662_ sky130_fd_sc_hd__mux2_2
XFILLER_0_166_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_511 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_15_596 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22204_ VGND VPWR _06589_ _06553_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_127_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23184_ VGND VPWR VGND VPWR _07079_ _03643_ _03642_ _03646_ _07011_ sky130_fd_sc_hd__a211o_2
XFILLER_0_28_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20396_ VGND VPWR _00966_ _05625_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_258_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_203_1112 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_24_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22135_ VPWR VGND _08933_ _06551_ _05385_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_30_577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_259_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22066_ VPWR VGND keymem.key_mem\[3\]\[95\] _06515_ _06405_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_255_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21017_ VGND VPWR VPWR VGND _05956_ _05066_ keymem.key_mem\[7\]\[116\] _05957_ sky130_fd_sc_hd__mux2_2
XFILLER_0_261_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_199_524 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_138_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25825_ VGND VPWR VPWR VGND clk _02318_ reset_n enc_block.block_w3_reg\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_177_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13770_ VGND VPWR VGND VPWR _09242_ enc_block.block_w2_reg\[24\] enc_block.sword_ctr_reg\[1\]
+ enc_block.sword_ctr_reg\[0\] sky130_fd_sc_hd__and3b_2
X_25756_ keymem.prev_key1_reg\[72\] clk _02249_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22968_ VGND VPWR VGND VPWR _02215_ _06948_ _06916_ keymem.prev_key1_reg\[38\] sky130_fd_sc_hd__o21a_2
XFILLER_0_74_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12721_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[55\] _08259_ _08268_ _08263_ _08269_
+ sky130_fd_sc_hd__o22a_2
X_24707_ VGND VPWR VPWR VGND clk _01200_ reset_n keymem.key_mem\[7\]\[60\] sky130_fd_sc_hd__dfrtp_2
X_21919_ VPWR VGND keymem.key_mem\[3\]\[26\] _06437_ _06427_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_179_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_70_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25687_ keymem.prev_key1_reg\[3\] clk _02180_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22899_ VGND VPWR VGND VPWR _11029_ _06890_ _11038_ _06905_ sky130_fd_sc_hd__a21o_2
XFILLER_0_35_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15440_ VGND VPWR VPWR VGND _10901_ _10735_ _10898_ _10899_ _10900_ sky130_fd_sc_hd__o31a_2
X_12652_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[49\] _07597_ keymem.key_mem\[7\]\[49\]
+ _07703_ _08206_ sky130_fd_sc_hd__a22o_2
X_24638_ VGND VPWR VPWR VGND clk _01131_ reset_n keymem.key_mem\[8\]\[119\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15371_ VGND VPWR _10832_ _10092_ _10833_ _10829_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_24569_ VGND VPWR VPWR VGND clk _01062_ reset_n keymem.key_mem\[8\]\[50\] sky130_fd_sc_hd__dfrtp_2
X_12583_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[42\] _07893_ _08143_ _08136_ _08144_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_0_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14322_ VGND VPWR _09792_ keymem.prev_key1_reg\[66\] _09791_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_17110_ VGND VPWR VPWR VGND _03220_ keylen _03226_ _03225_ _03224_ sky130_fd_sc_hd__o211a_2
X_18090_ VGND VPWR _04009_ enc_block.block_w0_reg\[26\] enc_block.block_w0_reg\[31\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1050 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_68_1167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_135_384 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17041_ VGND VPWR _00073_ _03163_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_149_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14253_ VPWR VGND VPWR VGND _09723_ _09638_ _09636_ key[129] _09544_ _09724_ sky130_fd_sc_hd__a221o_2
XFILLER_0_150_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_145_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_150_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13204_ VGND VPWR VGND VPWR _07793_ keymem.key_mem\[0\]\[103\] _08703_ _08699_ _08697_
+ _08704_ sky130_fd_sc_hd__o32a_2
XFILLER_0_81_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14184_ VGND VPWR VGND VPWR _09115_ _09097_ _09655_ _09077_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_106_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13135_ VGND VPWR enc_block.round_key\[96\] _08641_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18992_ VGND VPWR _04823_ _04753_ _04822_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_249_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1020 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13066_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[90\] _07685_ keymem.key_mem\[4\]\[90\]
+ _07636_ _08579_ sky130_fd_sc_hd__a22o_2
X_17943_ VGND VPWR VPWR VGND _03876_ key[233] keymem.prev_key1_reg\[105\] _03893_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_253_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12017_ VGND VPWR _07619_ _07618_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_246_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17874_ VGND VPWR VGND VPWR _03352_ keymem.prev_key1_reg\[83\] _03846_ _03818_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_217_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_40_1086 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19613_ VGND VPWR _00599_ _05209_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_178_1199 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16825_ VGND VPWR VGND VPWR _02967_ _02928_ _02927_ key[42] sky130_fd_sc_hd__o21a_2
XFILLER_0_205_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_156_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_878 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_136_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_215_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_117_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19544_ VGND VPWR _05173_ _05094_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_156_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16756_ VGND VPWR VPWR VGND _02884_ keymem.key_mem\[14\]\[35\] _02904_ _02905_ sky130_fd_sc_hd__mux2_2
X_13968_ VGND VPWR _09440_ _09439_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_92_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15707_ VGND VPWR VGND VPWR _11163_ enc_block.block_w2_reg\[18\] enc_block.sword_ctr_reg\[1\]
+ enc_block.sword_ctr_reg\[0\] sky130_fd_sc_hd__and3b_2
X_19475_ VGND VPWR VGND VPWR _05136_ keymem.key_mem_we _02894_ _05135_ _00534_ sky130_fd_sc_hd__a31o_2
X_12919_ VGND VPWR VGND VPWR _08447_ _07721_ keymem.key_mem\[14\]\[75\] _08444_ _08446_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_5_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13899_ VPWR VGND VGND VPWR _09371_ _09300_ _09246_ sky130_fd_sc_hd__nand2_2
X_16687_ VGND VPWR _00042_ _02840_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_9_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18426_ VPWR VGND VGND VPWR _04304_ _04314_ _03949_ sky130_fd_sc_hd__nor2_2
XFILLER_0_236_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_181_1_Left_448 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15638_ VGND VPWR VGND VPWR _11095_ _10189_ _11094_ _11092_ _11096_ sky130_fd_sc_hd__a31o_2
XFILLER_0_5_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_655 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18357_ _04251_ _04253_ _04008_ _04252_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_51_1182 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15569_ VGND VPWR VGND VPWR _09517_ _11026_ _11024_ _11025_ _11028_ sky130_fd_sc_hd__a31o_2
XFILLER_0_51_1193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_43_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17308_ VPWR VGND VPWR VGND _03403_ keymem.prev_key0_reg\[89\] sky130_fd_sc_hd__inv_2
X_18288_ VPWR VGND VPWR VGND _04191_ _03970_ _02394_ sky130_fd_sc_hd__or2_2
XFILLER_0_167_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_744 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17239_ VPWR VGND VPWR VGND _03341_ key[210] sky130_fd_sc_hd__inv_2
XFILLER_0_128_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_163_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20250_ VGND VPWR _00896_ _05549_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_25_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_204_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_163_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1565 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_243_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20181_ VGND VPWR VPWR VGND _05504_ _03555_ keymem.key_mem\[10\]\[110\] _05511_ sky130_fd_sc_hd__mux2_2
XFILLER_0_25_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_204_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_43_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23940_ VGND VPWR VPWR VGND clk _00433_ reset_n keymem.key_mem\[13\]\[61\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23871_ VGND VPWR VPWR VGND clk _00364_ reset_n enc_block.block_w2_reg\[24\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_174_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25610_ VGND VPWR VPWR VGND clk _02103_ reset_n keymem.key_mem\[0\]\[67\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_135_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22822_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[121\] _06860_ _06859_ _05077_ _02157_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_196_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_174_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_71_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_135_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25541_ VGND VPWR VPWR VGND clk _02034_ reset_n keymem.key_mem\[1\]\[126\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22753_ VGND VPWR VPWR VGND _06833_ keymem.key_mem\[0\]\[71\] _03252_ _06842_ sky130_fd_sc_hd__mux2_2
XFILLER_0_250_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_1093 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_920 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21704_ VGND VPWR _01578_ _06321_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_266_Right_135 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25472_ VGND VPWR VPWR VGND clk _01965_ reset_n keymem.key_mem\[1\]\[57\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_48_953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_66_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22684_ VGND VPWR VPWR VGND _06809_ keymem.key_mem\[0\]\[30\] _02839_ _06814_ sky130_fd_sc_hd__mux2_2
X_24423_ VGND VPWR VPWR VGND clk _00916_ reset_n keymem.key_mem\[9\]\[32\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_211_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21635_ VGND VPWR VPWR VGND _06275_ _02607_ keymem.key_mem\[4\]\[22\] _06285_ sky130_fd_sc_hd__mux2_2
XFILLER_0_19_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_474 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_945 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_198 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24354_ VGND VPWR VPWR VGND clk _00847_ reset_n keymem.key_mem\[10\]\[91\] sky130_fd_sc_hd__dfrtp_2
X_21566_ VGND VPWR _01514_ _06247_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23305_ VGND VPWR _07186_ enc_block.block_w2_reg\[1\] enc_block.block_w2_reg\[2\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_989 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_132_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20517_ VPWR VGND VGND VPWR _05676_ _05690_ keymem.key_mem\[8\]\[11\] sky130_fd_sc_hd__nor2_2
XFILLER_0_50_628 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24285_ VGND VPWR VPWR VGND clk _00778_ reset_n keymem.key_mem\[10\]\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_15_360 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21497_ VGND VPWR _01481_ _06211_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_144_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_181_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23236_ VPWR VGND VPWR VGND _07123_ block[3] _04837_ enc_block.block_w2_reg\[3\]
+ _04798_ _07124_ sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_164_2_Right_236 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20448_ VGND VPWR VPWR VGND _05649_ _03538_ keymem.key_mem\[9\]\[107\] _05653_ sky130_fd_sc_hd__mux2_2
XFILLER_0_142_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_28_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23167_ VGND VPWR _02294_ _07068_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20379_ VPWR VGND VGND VPWR _05617_ keymem.key_mem\[9\]\[74\] _05532_ sky130_fd_sc_hd__nand2_2
XFILLER_0_222_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22118_ VGND VPWR _01771_ _06542_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23098_ VGND VPWR _02268_ _07025_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_228_970 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14940_ enc_block.sword_ctr_reg\[1\] _10404_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[11\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_22049_ VGND VPWR _01738_ _06506_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_237_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14871_ VGND VPWR VGND VPWR _10172_ _10335_ _10336_ _09220_ _10332_ sky130_fd_sc_hd__nor4_2
XFILLER_0_255_1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_214_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16610_ VGND VPWR _00039_ _02766_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13822_ VGND VPWR _09294_ _09293_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_215_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25808_ keymem.prev_key1_reg\[124\] clk _02301_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_17590_ VPWR VGND VGND VPWR _03649_ _03240_ _02793_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13753_ VPWR VGND VGND VPWR _09222_ _09225_ _09067_ sky130_fd_sc_hd__nor2_2
XFILLER_0_74_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16541_ VPWR VGND VPWR VGND _02700_ keymem.prev_key0_reg\[121\] sky130_fd_sc_hd__inv_2
XFILLER_0_35_1133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25739_ keymem.prev_key1_reg\[55\] clk _02232_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_6_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12704_ VPWR VGND VPWR VGND _08252_ keymem.key_mem\[14\]\[54\] _08032_ keymem.key_mem\[11\]\[54\]
+ _07781_ _08253_ sky130_fd_sc_hd__a221o_2
X_19260_ VGND VPWR VPWR VGND _04993_ _05002_ keymem.key_mem\[13\]\[81\] _05003_ sky130_fd_sc_hd__mux2_2
X_16472_ VGND VPWR VGND VPWR _11352_ _11295_ _11275_ _11222_ _11252_ _02633_ sky130_fd_sc_hd__o32a_2
XFILLER_0_35_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13684_ VGND VPWR _09156_ _09135_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_6_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_233_Right_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18211_ VPWR VGND VGND VPWR _04120_ _04045_ _04119_ sky130_fd_sc_hd__nand2_2
X_15423_ VGND VPWR VGND VPWR _10883_ _10638_ _10884_ _10672_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_127_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12635_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[47\] _08145_ _08190_ _08186_ _08191_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_2_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19191_ VGND VPWR _04961_ _04879_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_249_1145 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_38_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1446 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18142_ VPWR VGND VGND VPWR _04057_ enc_block.block_w3_reg\[6\] _04056_ sky130_fd_sc_hd__nand2_2
X_15354_ _09827_ _10816_ _07386_ _09850_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_65_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12566_ VPWR VGND VPWR VGND _08127_ keymem.key_mem\[3\]\[41\] _07844_ keymem.key_mem\[12\]\[41\]
+ _07807_ _08128_ sky130_fd_sc_hd__a221o_2
XFILLER_0_31_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14305_ VPWR VGND VGND VPWR _09775_ _09773_ _09774_ sky130_fd_sc_hd__nand2_2
XFILLER_0_41_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18073_ VPWR VGND VPWR VGND _03994_ _03970_ _10666_ sky130_fd_sc_hd__or2_2
X_15285_ VGND VPWR VPWR VGND _09864_ keymem.key_mem\[14\]\[9\] _10747_ _10748_ sky130_fd_sc_hd__mux2_2
XFILLER_0_13_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12497_ VGND VPWR enc_block.round_key\[34\] _08065_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14236_ VGND VPWR VGND VPWR _09038_ _09707_ _09703_ _09706_ _09699_ sky130_fd_sc_hd__and4bb_2
X_17024_ VPWR VGND VPWR VGND _03148_ _10086_ _03145_ _03146_ _03147_ _10096_ sky130_fd_sc_hd__o311a_2
XFILLER_0_1_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_853 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_46_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14167_ VGND VPWR _09638_ _09637_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_238_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13118_ VPWR VGND VPWR VGND _08625_ keymem.key_mem\[6\]\[95\] _07739_ keymem.key_mem\[4\]\[95\]
+ _07914_ _08626_ sky130_fd_sc_hd__a221o_2
X_18975_ VGND VPWR _04808_ enc_block.block_w0_reg\[15\] _04807_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_14098_ VGND VPWR VGND VPWR _09391_ _09565_ _09569_ _09396_ sky130_fd_sc_hd__a21oi_2
X_17926_ VGND VPWR VPWR VGND _03874_ _03881_ keymem.prev_key0_reg\[99\] _03882_ sky130_fd_sc_hd__mux2_2
X_13049_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[88\] _07694_ keymem.key_mem\[11\]\[88\]
+ _07861_ _08564_ sky130_fd_sc_hd__a22o_2
XFILLER_0_186_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_147_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_480 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_56_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17857_ VGND VPWR _00218_ _03834_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16808_ VGND VPWR VGND VPWR _10379_ _10375_ _02952_ _02951_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_206_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_117_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17788_ _03675_ _03787_ _03106_ _03786_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_156_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19527_ VGND VPWR _05164_ _05092_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16739_ VGND VPWR VPWR VGND _09853_ _09854_ _09516_ _02889_ sky130_fd_sc_hd__or3_2
XFILLER_0_117_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19458_ VPWR VGND keymem.key_mem\[12\]\[27\] _05127_ _05116_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_18_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18409_ VPWR VGND _04300_ _04299_ enc_block.round_key\[127\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_88_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19389_ VPWR VGND keymem.key_mem_we _05087_ _03661_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_267_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21420_ VGND VPWR VPWR VGND _06162_ _03046_ keymem.key_mem\[5\]\[49\] _06171_ sky130_fd_sc_hd__mux2_2
XFILLER_0_71_252 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_44_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21351_ VGND VPWR VPWR VGND _06128_ _11446_ keymem.key_mem\[5\]\[16\] _06135_ sky130_fd_sc_hd__mux2_2
XFILLER_0_31_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1037 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20302_ VGND VPWR _00921_ _05576_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_128_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24070_ VGND VPWR VPWR VGND clk _00563_ reset_n keymem.key_mem\[12\]\[63\] sky130_fd_sc_hd__dfrtp_2
X_21282_ VGND VPWR VPWR VGND _06087_ _03573_ keymem.key_mem\[6\]\[113\] _06097_ sky130_fd_sc_hd__mux2_2
XFILLER_0_188_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_124_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23021_ VPWR VGND VPWR VGND _06980_ keymem.prev_key1_reg\[60\] _06926_ sky130_fd_sc_hd__or2_2
XFILLER_0_29_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20233_ VGND VPWR _00888_ _05540_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_13_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_756 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_228_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20164_ VGND VPWR VPWR VGND _05493_ _03506_ keymem.key_mem\[10\]\[102\] _05502_ sky130_fd_sc_hd__mux2_2
XFILLER_0_256_564 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_99_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24972_ VGND VPWR VPWR VGND clk _01465_ reset_n keymem.key_mem\[5\]\[69\] sky130_fd_sc_hd__dfrtp_2
X_20095_ VGND VPWR VPWR VGND _05457_ _03235_ keymem.key_mem\[10\]\[69\] _05466_ sky130_fd_sc_hd__mux2_2
X_23923_ VGND VPWR VPWR VGND clk _00416_ reset_n keymem.key_mem\[13\]\[44\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_1144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_97_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23854_ VGND VPWR VPWR VGND clk _00347_ reset_n enc_block.block_w2_reg\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_98_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_135_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1214 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_212_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22805_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[106\] _06858_ _06857_ _05045_ _02142_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_71_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23785_ VGND VPWR VPWR VGND clk _00278_ reset_n enc_block.block_w0_reg\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_75_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20997_ VGND VPWR _01246_ _05946_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_223_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22736_ VGND VPWR _06833_ _06778_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25524_ VGND VPWR VPWR VGND clk _02017_ reset_n keymem.key_mem\[1\]\[109\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_199 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25455_ VGND VPWR VPWR VGND clk _01948_ reset_n keymem.key_mem\[1\]\[40\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_94_388 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22667_ VGND VPWR VPWR VGND _06798_ keymem.key_mem\[0\]\[22\] _02608_ _06805_ sky130_fd_sc_hd__mux2_2
XFILLER_0_48_783 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_1030 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12420_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[28\] _07577_ keymem.key_mem\[4\]\[28\]
+ _07550_ _07995_ sky130_fd_sc_hd__a22o_2
X_24406_ VGND VPWR VPWR VGND clk _00899_ reset_n keymem.key_mem\[9\]\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_433 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21618_ VGND VPWR _01537_ _06276_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_30_1063 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_293 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25386_ VGND VPWR VPWR VGND clk _01879_ reset_n keymem.key_mem\[2\]\[99\] sky130_fd_sc_hd__dfrtp_2
X_22598_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[110\] _06775_ _06774_ _05054_ _02018_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_36_989 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_915 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24337_ VGND VPWR VPWR VGND clk _00830_ reset_n keymem.key_mem\[10\]\[74\] sky130_fd_sc_hd__dfrtp_2
X_12351_ VGND VPWR VGND VPWR _07933_ _07552_ keymem.key_mem\[4\]\[21\] _07930_ _07932_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_1_1484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21549_ VGND VPWR _01506_ _06238_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_35_488 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_691 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15070_ VPWR VGND VPWR VGND _10457_ _10445_ _10430_ _10419_ _10534_ sky130_fd_sc_hd__or4_2
X_12282_ VGND VPWR VGND VPWR _07869_ _07584_ keymem.key_mem\[14\]\[16\] _07866_ _07868_
+ sky130_fd_sc_hd__a211o_2
X_24268_ VGND VPWR VPWR VGND clk _00761_ reset_n keymem.key_mem\[10\]\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_205_1015 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_146_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1026 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14021_ VPWR VGND VGND VPWR _09397_ _09378_ _09493_ _09444_ _09416_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_82_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_165_2_Right_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23219_ VGND VPWR _07108_ enc_block.block_w0_reg\[18\] _07107_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_24199_ VGND VPWR VPWR VGND clk _00692_ reset_n keymem.key_mem\[11\]\[64\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_43_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18760_ VPWR VGND VPWR VGND _04614_ _04550_ _04612_ enc_block.block_w2_reg\[1\] _04602_
+ _00341_ sky130_fd_sc_hd__a221o_2
XFILLER_0_257_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15972_ VGND VPWR VGND VPWR _11428_ _11426_ _11221_ _11427_ _11365_ _11356_ sky130_fd_sc_hd__a32o_2
XFILLER_0_219_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17711_ VGND VPWR VGND VPWR _03740_ keymem.prev_key0_reg\[25\] _00166_ _03736_ sky130_fd_sc_hd__a21bo_2
X_14923_ VGND VPWR _10387_ _09021_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_257_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18691_ VGND VPWR _04552_ enc_block.block_w2_reg\[18\] enc_block.block_w0_reg\[3\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_984 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17642_ VGND VPWR _00147_ _03690_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_264_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14854_ VPWR VGND _10319_ keymem.prev_key1_reg\[39\] keymem.prev_key1_reg\[7\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_118_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13805_ VGND VPWR VGND VPWR _09277_ enc_block.block_w2_reg\[30\] enc_block.sword_ctr_reg\[1\]
+ enc_block.sword_ctr_reg\[0\] sky130_fd_sc_hd__and3b_2
XFILLER_0_114_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_453 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17573_ VGND VPWR _00134_ _03634_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_187_346 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14785_ VGND VPWR VGND VPWR _09357_ _09391_ _09363_ _09311_ _09373_ _10251_ sky130_fd_sc_hd__o32a_2
XFILLER_0_58_514 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11997_ VGND VPWR _07600_ _07599_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_54_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19312_ VPWR VGND keymem.key_mem_we _05035_ _03499_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16524_ _02682_ _02684_ _02681_ _02683_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_13736_ VPWR VGND VGND VPWR _09122_ _09208_ _09146_ sky130_fd_sc_hd__nor2_2
XFILLER_0_15_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_761 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19243_ VGND VPWR VPWR VGND _00447_ _04880_ _03286_ _08922_ _04991_ sky130_fd_sc_hd__o31ai_2
X_16455_ VPWR VGND VPWR VGND _02580_ _02615_ _02614_ _02576_ _02616_ sky130_fd_sc_hd__or4_2
X_13667_ VGND VPWR VPWR VGND _08963_ _08971_ _09009_ _09139_ sky130_fd_sc_hd__or3_2
XFILLER_0_229_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_945 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15406_ VGND VPWR _10867_ _10611_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12618_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[46\] _07760_ keymem.key_mem\[12\]\[46\]
+ _07722_ _08175_ sky130_fd_sc_hd__a22o_2
X_19174_ VPWR VGND keymem.key_mem_we _04950_ _03035_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13598_ VPWR VGND VGND VPWR _09067_ _09007_ _09070_ _09069_ _08999_ sky130_fd_sc_hd__o22ai_2
X_16386_ VPWR VGND VPWR VGND _02548_ _02497_ _02495_ key[149] _11043_ _02549_ sky130_fd_sc_hd__a221o_2
XFILLER_0_264_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1276 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18125_ VPWR VGND VGND VPWR _04042_ _04004_ _10185_ sky130_fd_sc_hd__nand2_2
X_15337_ VGND VPWR VGND VPWR _10628_ _10574_ _10565_ _10629_ _10799_ sky130_fd_sc_hd__o22a_2
XFILLER_0_5_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12549_ VGND VPWR VGND VPWR _08113_ _07712_ keymem.key_mem\[6\]\[39\] _08110_ _08112_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_13_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_108_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_262_1131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_101_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_125_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18056_ VGND VPWR _03977_ _03947_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_164_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15268_ VGND VPWR _10731_ keymem.prev_key0_reg\[105\] _10730_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_125_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17007_ VPWR VGND _03132_ _02751_ _02750_ VPWR VGND sky130_fd_sc_hd__xor2_2
X_14219_ VGND VPWR VGND VPWR _09102_ _09173_ _09077_ _09108_ _09230_ _09690_ sky130_fd_sc_hd__o32a_2
XFILLER_0_50_981 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_61_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15199_ VGND VPWR VPWR VGND _09864_ keymem.key_mem\[14\]\[8\] _10662_ _10663_ sky130_fd_sc_hd__mux2_2
XFILLER_0_111_357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_201_1446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_201_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18958_ VGND VPWR _04793_ _04791_ _04792_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_236_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17909_ VGND VPWR VGND VPWR _03792_ _02830_ _03727_ _03859_ _03870_ _03794_ sky130_fd_sc_hd__a2111o_2
X_18889_ VGND VPWR VGND VPWR _04729_ _04728_ _04731_ _04727_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_222_910 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20920_ VGND VPWR VPWR VGND _05880_ _04983_ keymem.key_mem\[7\]\[70\] _05906_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_125_1_Left_392 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_90_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_95_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20851_ VGND VPWR VGND VPWR _05869_ keymem.key_mem_we _02924_ _05864_ _01177_ sky130_fd_sc_hd__a31o_2
XFILLER_0_132_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23570_ VGND VPWR VPWR VGND clk _00071_ reset_n keymem.key_mem\[14\]\[59\] sky130_fd_sc_hd__dfrtp_2
X_20782_ VPWR VGND keymem.key_mem\[7\]\[6\] _05832_ _05830_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_212_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22521_ VGND VPWR VPWR VGND _06739_ keymem.key_mem\[1\]\[61\] _03162_ _06748_ sky130_fd_sc_hd__mux2_2
XFILLER_0_64_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_130_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25240_ VGND VPWR VPWR VGND clk _01733_ reset_n keymem.key_mem\[3\]\[81\] sky130_fd_sc_hd__dfrtp_2
X_22452_ VGND VPWR VPWR VGND _06715_ keymem.key_mem\[1\]\[20\] _02480_ _06720_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_444 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_161_213 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_267_1086 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21403_ VGND VPWR _06162_ _06116_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_228_1037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25171_ VGND VPWR VPWR VGND clk _01664_ reset_n keymem.key_mem\[3\]\[12\] sky130_fd_sc_hd__dfrtp_2
X_22383_ VGND VPWR VPWR VGND _06680_ _03592_ keymem.key_mem\[2\]\[116\] _06683_ sky130_fd_sc_hd__mux2_2
XFILLER_0_161_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24122_ VGND VPWR VPWR VGND clk _00615_ reset_n keymem.key_mem\[12\]\[115\] sky130_fd_sc_hd__dfrtp_2
X_21334_ VGND VPWR VPWR VGND _06117_ _10661_ keymem.key_mem\[5\]\[8\] _06126_ sky130_fd_sc_hd__mux2_2
XFILLER_0_128_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_382 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_335 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24053_ VGND VPWR VPWR VGND clk _00546_ reset_n keymem.key_mem\[12\]\[46\] sky130_fd_sc_hd__dfrtp_2
X_21265_ VGND VPWR _01372_ _06088_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23004_ VGND VPWR VPWR VGND _06960_ _03081_ keymem.prev_key1_reg\[53\] _06970_ sky130_fd_sc_hd__mux2_2
XFILLER_0_102_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20216_ VGND VPWR VPWR VGND _05388_ _03668_ keymem.key_mem\[10\]\[127\] _05529_ sky130_fd_sc_hd__mux2_2
XFILLER_0_12_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_60_1045 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_99_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21196_ VGND VPWR _06052_ _05970_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_60_1067 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_501 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_218_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20147_ VGND VPWR _05493_ _05387_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_229_597 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_217_737 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20078_ VGND VPWR _05457_ _05387_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24955_ VGND VPWR VPWR VGND clk _01448_ reset_n keymem.key_mem\[5\]\[52\] sky130_fd_sc_hd__dfrtp_2
X_11920_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[31\] dec_new_block\[127\]
+ _07524_ sky130_fd_sc_hd__mux2_2
X_23906_ VGND VPWR VPWR VGND clk _00399_ reset_n keymem.key_mem\[13\]\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_197_600 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24886_ VGND VPWR VPWR VGND clk _01379_ reset_n keymem.key_mem\[6\]\[111\] sky130_fd_sc_hd__dfrtp_2
X_11851_ VGND VPWR result[92] _07489_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23837_ VGND VPWR VPWR VGND clk _00330_ reset_n enc_block.block_w1_reg\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_213_987 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_212_486 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14570_ VGND VPWR VGND VPWR _09350_ _09358_ _09305_ _09576_ _10038_ sky130_fd_sc_hd__o22a_2
XFILLER_0_36_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11782_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[26\] dec_new_block\[58\]
+ _07455_ sky130_fd_sc_hd__mux2_2
X_23768_ keymem.prev_key0_reg\[124\] clk _00265_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_3_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13521_ enc_block.sword_ctr_reg\[1\] _08993_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[4\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_25507_ VGND VPWR VPWR VGND clk _02000_ reset_n keymem.key_mem\[1\]\[92\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22719_ VGND VPWR VPWR VGND _06822_ keymem.key_mem\[0\]\[54\] _03091_ _06825_ sky130_fd_sc_hd__mux2_2
X_23699_ keymem.prev_key0_reg\[55\] clk _00196_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_211_1074 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16240_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[51\] keymem.prev_key1_reg\[19\]
+ _02404_ _02405_ sky130_fd_sc_hd__a21o_2
X_13452_ VPWR VGND VPWR VGND _08924_ keymem.round_ctr_reg\[0\] keymem.round_ctr_reg\[1\]
+ sky130_fd_sc_hd__or2_2
X_25438_ VGND VPWR VPWR VGND clk _01931_ reset_n keymem.key_mem\[1\]\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12403_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[26\] _07608_ keymem.key_mem\[14\]\[26\]
+ _07582_ _07980_ sky130_fd_sc_hd__a22o_2
X_16171_ VPWR VGND VPWR VGND _11561_ _02337_ _11624_ _11622_ sky130_fd_sc_hd__or3b_2
X_25369_ VGND VPWR VPWR VGND clk _01862_ reset_n keymem.key_mem\[2\]\[82\] sky130_fd_sc_hd__dfrtp_2
X_13383_ VGND VPWR VGND VPWR _08865_ _08096_ keymem.key_mem\[5\]\[121\] _08862_ _08864_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_23_414 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15122_ VPWR VGND VPWR VGND _10424_ _10445_ _10430_ _10419_ _10586_ sky130_fd_sc_hd__or4_2
X_12334_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[20\] _07845_ keymem.key_mem\[14\]\[20\]
+ _07782_ _07917_ sky130_fd_sc_hd__a22o_2
XFILLER_0_107_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15053_ VPWR VGND VGND VPWR _10513_ _10515_ _10516_ _10517_ sky130_fd_sc_hd__nor3_2
X_19930_ VGND VPWR _00748_ _05377_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_50_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12265_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[15\] _07619_ keymem.key_mem\[12\]\[15\]
+ _07722_ _07853_ sky130_fd_sc_hd__a22o_2
XFILLER_0_107_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14004_ VGND VPWR _09476_ _09434_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_166_2_Right_238 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_142_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19861_ VGND VPWR _00715_ _05341_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12196_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[10\] _07695_ keymem.key_mem\[12\]\[10\]
+ _07788_ _07789_ sky130_fd_sc_hd__a22o_2
XFILLER_0_222_1181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18812_ VPWR VGND VPWR VGND _04661_ block[38] _04576_ enc_block.block_w1_reg\[6\]
+ _04543_ _04662_ sky130_fd_sc_hd__a221o_2
XFILLER_0_128_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_821 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_190_1_Left_457 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19792_ VGND VPWR _00682_ _05305_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_207_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_78_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18743_ VPWR VGND VGND VPWR _04305_ _04599_ _03948_ sky130_fd_sc_hd__nor2_2
X_15955_ VGND VPWR VGND VPWR _11218_ _11316_ _11411_ _11238_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_120_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_263_887 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_257_1277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_262_386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14906_ VGND VPWR _00019_ _10370_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18674_ VGND VPWR _04537_ _04320_ _04471_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15886_ VGND VPWR VGND VPWR _11333_ _11323_ _11335_ _11337_ _11342_ _11341_ sky130_fd_sc_hd__a2111o_2
X_17625_ VGND VPWR _00142_ _03678_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_118_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14837_ VGND VPWR VGND VPWR _09410_ _09294_ _10302_ _09476_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_77_119 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_15_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17556_ VPWR VGND VPWR VGND _03619_ _03616_ _03615_ key[248] _08929_ _03620_ sky130_fd_sc_hd__a221o_2
X_14768_ VPWR VGND VPWR VGND _10234_ _09435_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_128_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16507_ VPWR VGND VGND VPWR keymem.prev_key0_reg\[120\] _02666_ _07387_ _02664_ _02665_
+ _02667_ sky130_fd_sc_hd__a311o_2
X_13719_ _09190_ _09191_ _09189_ _09188_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_17487_ VPWR VGND VPWR VGND _03559_ _03557_ _03020_ key[239] _03527_ _03560_ sky130_fd_sc_hd__a221o_2
X_14699_ VPWR VGND VGND VPWR _10166_ _10165_ _10163_ _09806_ _09178_ _09095_ sky130_fd_sc_hd__o2111a_2
XFILLER_0_89_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19226_ VGND VPWR VPWR VGND _00440_ _04880_ _03226_ _08922_ _04981_ sky130_fd_sc_hd__o31ai_2
X_16438_ _02597_ _02600_ keymem.prev_key1_reg\[86\] _02598_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_89_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19157_ VPWR VGND keymem.key_mem_we _04939_ _02972_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_143_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16369_ VGND VPWR VGND VPWR _11327_ _11352_ _02532_ _11465_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_27_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18108_ VGND VPWR _04026_ _04023_ _04025_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_19088_ VGND VPWR VGND VPWR _04898_ keymem.key_mem_we _11040_ _04896_ _00385_ sky130_fd_sc_hd__a31o_2
XFILLER_0_48_1165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_125_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_615 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18039_ VGND VPWR _03961_ enc_block.block_w2_reg\[8\] enc_block.block_w1_reg\[16\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_257_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_199_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21050_ VGND VPWR _01270_ _05975_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_26_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_396 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_10_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20001_ VGND VPWR VPWR VGND _05413_ _02689_ keymem.key_mem\[10\]\[24\] _05417_ sky130_fd_sc_hd__mux2_2
XFILLER_0_226_523 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_94_52 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_718 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_226_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_158_1153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21952_ VGND VPWR VPWR VGND _06449_ _04937_ keymem.key_mem\[3\]\[41\] _06455_ sky130_fd_sc_hd__mux2_2
X_24740_ VGND VPWR VPWR VGND clk _01233_ reset_n keymem.key_mem\[7\]\[93\] sky130_fd_sc_hd__dfrtp_2
X_20903_ VPWR VGND keymem.key_mem\[7\]\[62\] _05897_ _05886_ VPWR VGND sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_128_2_Right_200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24671_ VGND VPWR VPWR VGND clk _01164_ reset_n keymem.key_mem\[7\]\[24\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_136_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21883_ VGND VPWR VGND VPWR _06417_ keymem.key_mem_we _10747_ _06404_ _01661_ sky130_fd_sc_hd__a31o_2
XFILLER_0_33_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1085 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23622_ VGND VPWR VPWR VGND clk _00123_ reset_n keymem.key_mem\[14\]\[111\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_166_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20834_ VPWR VGND keymem.key_mem\[7\]\[30\] _05860_ _05856_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_37_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_76_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_76_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_193_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_37_517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23553_ VGND VPWR VPWR VGND clk _00054_ reset_n keymem.key_mem\[14\]\[42\] sky130_fd_sc_hd__dfrtp_2
X_20765_ VGND VPWR _05821_ _05820_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_9_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22504_ VGND VPWR _01959_ _06740_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_247_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23484_ VPWR VGND VGND VPWR _07345_ _07346_ _04382_ sky130_fd_sc_hd__nor2_2
XFILLER_0_91_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_68_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20696_ VGND VPWR VPWR VGND _05783_ _03466_ keymem.key_mem\[8\]\[96\] _05784_ sky130_fd_sc_hd__mux2_2
XFILLER_0_45_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25223_ VGND VPWR VPWR VGND clk _01716_ reset_n keymem.key_mem\[3\]\[64\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_247_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22435_ VGND VPWR VPWR VGND _06702_ keymem.key_mem\[1\]\[12\] _10977_ _06711_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25154_ VGND VPWR VPWR VGND clk _01647_ reset_n keymem.key_mem\[4\]\[123\] sky130_fd_sc_hd__dfrtp_2
X_22366_ VGND VPWR VPWR VGND _06669_ _03543_ keymem.key_mem\[2\]\[108\] _06674_ sky130_fd_sc_hd__mux2_2
XFILLER_0_21_929 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_108_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24105_ VGND VPWR VPWR VGND clk _00598_ reset_n keymem.key_mem\[12\]\[98\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21317_ VGND VPWR _06117_ _06116_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25085_ VGND VPWR VPWR VGND clk _01578_ reset_n keymem.key_mem\[4\]\[54\] sky130_fd_sc_hd__dfrtp_2
X_22297_ VPWR VGND VGND VPWR _06638_ keymem.key_mem\[2\]\[75\] _06567_ sky130_fd_sc_hd__nand2_2
XFILLER_0_44_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_248_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12050_ VGND VPWR _07650_ _07649_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24036_ VGND VPWR VPWR VGND clk _00529_ reset_n keymem.key_mem\[12\]\[29\] sky130_fd_sc_hd__dfrtp_2
X_21248_ VGND VPWR _01364_ _06079_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_236_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_178_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21179_ VGND VPWR _01331_ _06043_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_90_2_Right_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_258_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15740_ VPWR VGND VPWR VGND _11196_ enc_block.block_w0_reg\[20\] _08995_ sky130_fd_sc_hd__or2_2
XFILLER_0_245_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24938_ VGND VPWR VPWR VGND clk _01431_ reset_n keymem.key_mem\[5\]\[35\] sky130_fd_sc_hd__dfrtp_2
X_12952_ VGND VPWR enc_block.round_key\[78\] _08476_ VPWR VGND sky130_fd_sc_hd__buf_1
X_11903_ VGND VPWR result[118] _07515_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15671_ VGND VPWR VGND VPWR _10574_ _10575_ _10629_ _10478_ _10580_ _11128_ sky130_fd_sc_hd__o32a_2
XFILLER_0_169_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_73_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24869_ VGND VPWR VPWR VGND clk _01362_ reset_n keymem.key_mem\[6\]\[94\] sky130_fd_sc_hd__dfrtp_2
X_12883_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[72\] _07759_ keymem.key_mem\[9\]\[72\]
+ _07612_ _08414_ sky130_fd_sc_hd__a22o_2
XFILLER_0_115_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17410_ VGND VPWR _00112_ _03493_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14622_ VGND VPWR _10090_ keymem.prev_key1_reg\[4\] keymem.prev_key1_reg\[36\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
X_11834_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[20\] dec_new_block\[84\]
+ _07481_ sky130_fd_sc_hd__mux2_2
X_18390_ VPWR VGND VGND VPWR _04283_ _04004_ _10141_ sky130_fd_sc_hd__nand2_2
XFILLER_0_240_592 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_197_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_327 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_90_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_201_979 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_28_517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_67_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_200_467 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17341_ VGND VPWR VGND VPWR keylen _03433_ _03432_ _10371_ _02779_ _02780_ sky130_fd_sc_hd__a311oi_2
X_11765_ VGND VPWR result[49] _07446_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14553_ VGND VPWR VGND VPWR _09146_ _09138_ _10021_ _09109_ sky130_fd_sc_hd__a21oi_2
X_13504_ VPWR VGND VPWR VGND _08976_ enc_block.block_w0_reg\[7\] _08952_ sky130_fd_sc_hd__or2_2
X_17272_ VGND VPWR VPWR VGND _02488_ _02489_ _09868_ _03371_ sky130_fd_sc_hd__or3_2
XFILLER_0_265_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11696_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[15\] dec_new_block\[15\]
+ _07412_ sky130_fd_sc_hd__mux2_2
X_14484_ VGND VPWR VGND VPWR _09953_ _09687_ _09103_ _09067_ _09211_ _09952_ sky130_fd_sc_hd__o221ai_2
X_19011_ VPWR VGND VGND VPWR _04840_ _04625_ _04839_ sky130_fd_sc_hd__nand2_2
XFILLER_0_165_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16223_ VGND VPWR VGND VPWR _11392_ _11434_ _02385_ _02386_ _02388_ _02387_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_64_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13435_ VGND VPWR enc_block.round_key\[126\] _08911_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_10_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_723 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16154_ VPWR VGND VPWR VGND _11602_ _11607_ _11608_ _11595_ _11600_ sky130_fd_sc_hd__or4b_2
X_13366_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[120\] _08137_ keymem.key_mem\[9\]\[120\]
+ _07717_ _08849_ sky130_fd_sc_hd__a22o_2
XFILLER_0_10_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1232 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15105_ VGND VPWR _10569_ _10568_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_84_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12317_ VGND VPWR _07901_ _07714_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16085_ VPWR VGND VPWR VGND _11540_ keymem.prev_key0_reg\[17\] sky130_fd_sc_hd__inv_2
X_13297_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[113\] _07872_ keymem.key_mem\[11\]\[113\]
+ _07599_ _08787_ sky130_fd_sc_hd__a22o_2
XFILLER_0_267_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15036_ VGND VPWR _10500_ _10483_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12248_ VGND VPWR VGND VPWR _07542_ keymem.key_mem\[8\]\[14\] _07833_ _07836_ _07837_
+ _07574_ sky130_fd_sc_hd__a2111o_2
X_19913_ VGND VPWR _00740_ _05368_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_20_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_43_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_489 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_202_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_167_2_Right_239 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19844_ VGND VPWR _00707_ _05332_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12179_ VPWR VGND VPWR VGND _07772_ keymem.key_mem\[3\]\[9\] _07603_ keymem.key_mem\[6\]\[9\]
+ _07771_ _07773_ sky130_fd_sc_hd__a221o_2
XFILLER_0_120_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19775_ VGND VPWR _00674_ _05296_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16987_ _02712_ _03114_ keymem.prev_key1_reg\[57\] _02713_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_155_1304 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18726_ VPWR VGND VPWR VGND _04583_ _04550_ _04582_ enc_block.block_w1_reg\[30\]
+ _04328_ _00338_ sky130_fd_sc_hd__a221o_2
XFILLER_0_266_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15938_ VPWR VGND VPWR VGND _11393_ _11392_ _11390_ _11389_ _11290_ _11394_ sky130_fd_sc_hd__a221o_2
XFILLER_0_155_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1386 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_91_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_155_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18657_ VPWR VGND _04522_ _04372_ enc_block.block_w3_reg\[15\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15869_ VGND VPWR _11325_ _11324_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_91_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17608_ VPWR VGND VGND VPWR _03665_ _02852_ _02853_ sky130_fd_sc_hd__nand2_2
XFILLER_0_231_1236 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18588_ VPWR VGND VPWR VGND _04460_ _04459_ _04458_ enc_block.block_w1_reg\[15\]
+ _04424_ _00323_ sky130_fd_sc_hd__a221o_2
XFILLER_0_58_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17539_ VGND VPWR VGND VPWR _03604_ _10322_ _02597_ _02598_ _03605_ sky130_fd_sc_hd__a31o_2
XFILLER_0_73_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_104_61 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20550_ VGND VPWR _01038_ _05707_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_13_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_433 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_27_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19209_ VGND VPWR VGND VPWR _04971_ keymem.key_mem_we _03162_ _04968_ _00433_ sky130_fd_sc_hd__a31o_2
XFILLER_0_6_455 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_723 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20481_ VGND VPWR VPWR VGND _05660_ _03640_ keymem.key_mem\[9\]\[123\] _05670_ sky130_fd_sc_hd__mux2_2
XFILLER_0_7_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_211 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22220_ VGND VPWR _01818_ _06597_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_162_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_778 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_89_74 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_73_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22151_ VGND VPWR VPWR VGND _06554_ _10283_ keymem.key_mem\[2\]\[6\] _06561_ sky130_fd_sc_hd__mux2_2
XFILLER_0_30_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21102_ VGND VPWR VPWR VGND _05996_ _02764_ keymem.key_mem\[6\]\[27\] _06003_ sky130_fd_sc_hd__mux2_2
X_22082_ VGND VPWR _01754_ _06523_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_196_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_450 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21033_ VGND VPWR VPWR VGND _05956_ _05083_ keymem.key_mem\[7\]\[124\] _05965_ sky130_fd_sc_hd__mux2_2
XFILLER_0_201_1073 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25841_ VGND VPWR VPWR VGND clk _02334_ reset_n enc_block.block_w3_reg\[29\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_242_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_260_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22984_ VGND VPWR VGND VPWR _06958_ _03001_ _03000_ _03005_ _06951_ sky130_fd_sc_hd__a211o_2
X_25772_ keymem.prev_key1_reg\[88\] clk _02265_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_173_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24723_ VGND VPWR VPWR VGND clk _01216_ reset_n keymem.key_mem\[7\]\[76\] sky130_fd_sc_hd__dfrtp_2
X_21935_ VGND VPWR _01685_ _06445_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_215_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_2_Right_201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_171_1161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24654_ VGND VPWR VPWR VGND clk _01147_ reset_n keymem.key_mem\[7\]\[7\] sky130_fd_sc_hd__dfrtp_2
X_21866_ VGND VPWR VGND VPWR _06408_ keymem.key_mem_we _09725_ _06404_ _01653_ sky130_fd_sc_hd__a31o_2
XFILLER_0_132_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23605_ VGND VPWR VPWR VGND clk _00106_ reset_n keymem.key_mem\[14\]\[94\] sky130_fd_sc_hd__dfrtp_2
X_20817_ VPWR VGND keymem.key_mem\[7\]\[22\] _05851_ _05844_ VPWR VGND sky130_fd_sc_hd__and2_2
X_24585_ VGND VPWR VPWR VGND clk _01078_ reset_n keymem.key_mem\[8\]\[66\] sky130_fd_sc_hd__dfrtp_2
X_21797_ VGND VPWR VPWR VGND _06366_ _03485_ keymem.key_mem\[4\]\[99\] _06370_ sky130_fd_sc_hd__mux2_2
XFILLER_0_231_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23536_ VGND VPWR VPWR VGND clk _00037_ reset_n keymem.key_mem\[14\]\[25\] sky130_fd_sc_hd__dfrtp_2
X_20748_ VGND VPWR VPWR VGND _05805_ _03627_ keymem.key_mem\[8\]\[121\] _05811_ sky130_fd_sc_hd__mux2_2
XFILLER_0_110_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_147_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_52_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23467_ _07329_ _07331_ _03981_ _07330_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_110_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20679_ VGND VPWR VPWR VGND _05772_ _03401_ keymem.key_mem\[8\]\[88\] _05775_ sky130_fd_sc_hd__mux2_2
XFILLER_0_184_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13220_ VGND VPWR VGND VPWR _07593_ keymem.key_mem\[9\]\[105\] _08715_ _08717_ _08718_
+ _08599_ sky130_fd_sc_hd__a2111o_2
X_25206_ VGND VPWR VPWR VGND clk _01699_ reset_n keymem.key_mem\[3\]\[47\] sky130_fd_sc_hd__dfrtp_2
X_22418_ VGND VPWR _06702_ _06701_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_61_862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_162_385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23398_ VPWR VGND VPWR VGND block[19] _03979_ enc_block.block_w0_reg\[19\] _03977_
+ _07270_ sky130_fd_sc_hd__a22o_2
XFILLER_0_180_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_260_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13151_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[98\] _07651_ keymem.key_mem\[12\]\[98\]
+ _07787_ _08656_ sky130_fd_sc_hd__a22o_2
X_22349_ VGND VPWR VPWR VGND _06658_ _03492_ keymem.key_mem\[2\]\[100\] _06665_ sky130_fd_sc_hd__mux2_2
X_25137_ VGND VPWR VPWR VGND clk _01630_ reset_n keymem.key_mem\[4\]\[106\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_249_434 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_260_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1416 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12102_ VPWR VGND VPWR VGND _07699_ keymem.key_mem\[6\]\[5\] _07657_ keymem.key_mem\[2\]\[5\]
+ _07698_ _07700_ sky130_fd_sc_hd__a221o_2
X_13082_ VGND VPWR VGND VPWR _08594_ _07648_ keymem.key_mem\[2\]\[91\] _08591_ _08593_
+ sky130_fd_sc_hd__a211o_2
X_25068_ VGND VPWR VPWR VGND clk _01561_ reset_n keymem.key_mem\[4\]\[37\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_178_1304 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16910_ VGND VPWR VPWR VGND _03042_ _03039_ _03045_ _02496_ _03044_ sky130_fd_sc_hd__o211a_2
X_24019_ VGND VPWR VPWR VGND clk _00512_ reset_n keymem.key_mem\[12\]\[12\] sky130_fd_sc_hd__dfrtp_2
X_12033_ VPWR VGND VPWR VGND _07633_ keymem.key_mem\[14\]\[2\] _07632_ keymem.key_mem\[11\]\[2\]
+ _07631_ _07634_ sky130_fd_sc_hd__a221o_2
X_17890_ VGND VPWR VGND VPWR _03737_ keymem.prev_key1_reg\[88\] _03857_ _03738_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16841_ VPWR VGND key[171] _02982_ _09522_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_121_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_244_150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_233_824 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_91_2_Right_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_260_621 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_233_835 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_189_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19560_ VGND VPWR _00574_ _05181_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_191_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16772_ VPWR VGND VGND VPWR _10187_ _02919_ _10735_ sky130_fd_sc_hd__nor2_2
XFILLER_0_254_1236 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13984_ VGND VPWR _09456_ _09293_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18511_ VGND VPWR _04391_ _04062_ _00315_ _04317_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_15723_ VGND VPWR VGND VPWR _11179_ _11178_ _11177_ keymem.prev_key1_reg\[17\] _10402_
+ _09002_ sky130_fd_sc_hd__a32o_2
XFILLER_0_260_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12935_ VPWR VGND VPWR VGND _08460_ keymem.key_mem\[10\]\[77\] _07562_ keymem.key_mem\[4\]\[77\]
+ _08077_ _08461_ sky130_fd_sc_hd__a221o_2
X_19491_ VGND VPWR VPWR VGND _05138_ _04939_ keymem.key_mem\[12\]\[42\] _05145_ sky130_fd_sc_hd__mux2_2
XFILLER_0_125_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18442_ VPWR VGND VGND VPWR _04328_ _04329_ _03994_ sky130_fd_sc_hd__nor2_2
X_15654_ VGND VPWR _11111_ keymem.prev_key0_reg\[15\] _11110_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_12866_ VGND VPWR VGND VPWR _07835_ keymem.key_mem\[13\]\[70\] _08396_ _08398_ _08399_
+ _08243_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_200_220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_765 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14605_ VPWR VGND VPWR VGND _09590_ _09736_ _09604_ _09556_ _10073_ sky130_fd_sc_hd__or4_2
XFILLER_0_205_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11817_ VGND VPWR result[75] _07472_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18373_ VGND VPWR _04267_ _03976_ _00301_ _04258_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_200_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15585_ VGND VPWR _11043_ _09543_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12797_ VPWR VGND VPWR VGND keymem.key_mem\[6\]\[63\] _07760_ keymem.key_mem\[2\]\[63\]
+ _07816_ _08337_ sky130_fd_sc_hd__a22o_2
XFILLER_0_28_336 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_141_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17324_ VGND VPWR _03418_ _03417_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14536_ VGND VPWR VGND VPWR _09222_ _09160_ _09167_ _09116_ _10004_ sky130_fd_sc_hd__o22a_2
XFILLER_0_172_116 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11748_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[9\] dec_new_block\[41\]
+ _07438_ sky130_fd_sc_hd__mux2_2
XFILLER_0_56_689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17255_ VGND VPWR _03356_ _03355_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14467_ VPWR VGND VGND VPWR _09019_ _09936_ _09149_ sky130_fd_sc_hd__nor2_2
X_11679_ VGND VPWR result[6] _07403_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16206_ VPWR VGND VPWR VGND _02368_ _02370_ _02371_ _11416_ _11597_ sky130_fd_sc_hd__or4b_2
XFILLER_0_10_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13418_ VPWR VGND VPWR VGND _08895_ keymem.key_mem\[5\]\[125\] _07683_ keymem.key_mem\[9\]\[125\]
+ _07738_ _08896_ sky130_fd_sc_hd__a221o_2
XFILLER_0_148_1163 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_261_1229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17186_ key[204] _03294_ keylen _10325_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_14398_ VGND VPWR _09867_ keymem.prev_key1_reg\[3\] keymem.prev_key1_reg\[35\] VPWR
+ VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_226_1349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_180_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_49_1282 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16137_ VGND VPWR VGND VPWR _11469_ _11473_ _11591_ _11460_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_109_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13349_ VPWR VGND VPWR VGND keymem.key_mem\[12\]\[118\] _07787_ keymem.key_mem\[2\]\[118\]
+ _07697_ _08834_ sky130_fd_sc_hd__a22o_2
XFILLER_0_11_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_84_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_102_2_Left_573 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16068_ VGND VPWR VGND VPWR _11523_ _11392_ _11390_ _11368_ _11366_ sky130_fd_sc_hd__a211o_2
XFILLER_0_267_275 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_196_1404 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15019_ VGND VPWR _10483_ _10447_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_227_139 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_202_1382 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19827_ VGND VPWR _00699_ _05323_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_237_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_235_172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_247_Right_116 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_263_492 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19758_ VGND VPWR _00666_ _05287_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_223_345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_155_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18709_ VPWR VGND VPWR VGND _04568_ _04550_ _04567_ enc_block.block_w1_reg\[28\]
+ _04328_ _00336_ sky130_fd_sc_hd__a221o_2
X_19689_ VGND VPWR _00633_ _05251_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21720_ VGND VPWR _01586_ _06329_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_204_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_56_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_86 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21651_ VGND VPWR _01553_ _06293_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_46_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20602_ VGND VPWR _01063_ _05734_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24370_ VGND VPWR VPWR VGND clk _00863_ reset_n keymem.key_mem\[10\]\[107\] sky130_fd_sc_hd__dfrtp_2
X_21582_ VGND VPWR _01522_ _06255_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_129_382 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_35_829 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_129_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23321_ VGND VPWR _07201_ enc_block.round_key\[11\] _07200_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_248_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20533_ VGND VPWR _01030_ _05698_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23252_ VGND VPWR VPWR VGND _07093_ enc_block.block_w3_reg\[4\] _07138_ _07139_ sky130_fd_sc_hd__mux2_2
XFILLER_0_166_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20464_ VGND VPWR _00998_ _05661_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_171_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22203_ VGND VPWR _01810_ _06588_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23183_ VGND VPWR _02300_ _07078_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20395_ VGND VPWR VPWR VGND _05614_ _03347_ keymem.key_mem\[9\]\[82\] _05625_ sky130_fd_sc_hd__mux2_2
XFILLER_0_63_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22134_ VGND VPWR _01779_ _06550_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_144_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22065_ VGND VPWR _01746_ _06514_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_262_919 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21016_ VGND VPWR _05956_ _05819_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_227_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_103_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25824_ VGND VPWR VPWR VGND clk _02317_ reset_n enc_block.block_w3_reg\[12\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_173_1245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_241_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25755_ keymem.prev_key1_reg\[71\] clk _02248_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_69_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22967_ VGND VPWR VGND VPWR _06948_ _02929_ _02926_ _02933_ _06892_ sky130_fd_sc_hd__a211o_2
XFILLER_0_138_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_70_1206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24706_ VGND VPWR VPWR VGND clk _01199_ reset_n keymem.key_mem\[7\]\[59\] sky130_fd_sc_hd__dfrtp_2
X_12720_ VGND VPWR VGND VPWR _08268_ _08008_ keymem.key_mem\[2\]\[55\] _08264_ _08267_
+ sky130_fd_sc_hd__a211o_2
XPHY_EDGE_ROW_178_2_Left_649 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_69_258 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21918_ VGND VPWR VGND VPWR _06436_ keymem.key_mem_we _02721_ _06432_ _01677_ sky130_fd_sc_hd__a31o_2
X_25686_ keymem.prev_key1_reg\[2\] clk _02179_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22898_ VGND VPWR _02189_ _06904_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_70_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12651_ VGND VPWR VGND VPWR _07786_ keymem.key_mem\[10\]\[49\] _08202_ _08204_ _08205_
+ _08069_ sky130_fd_sc_hd__a2111o_2
X_24637_ VGND VPWR VPWR VGND clk _01130_ reset_n keymem.key_mem\[8\]\[118\] sky130_fd_sc_hd__dfrtp_2
X_21849_ VGND VPWR VPWR VGND _06388_ _03647_ keymem.key_mem\[4\]\[124\] _06397_ sky130_fd_sc_hd__mux2_2
XFILLER_0_37_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12582_ VGND VPWR VGND VPWR _08096_ keymem.key_mem\[5\]\[42\] _08138_ _08140_ _08143_
+ _08142_ sky130_fd_sc_hd__a2111o_2
X_15370_ VGND VPWR VGND VPWR _10832_ _10831_ _10830_ _09522_ sky130_fd_sc_hd__o21a_2
X_24568_ VGND VPWR VPWR VGND clk _01061_ reset_n keymem.key_mem\[8\]\[49\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_1313 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14321_ VGND VPWR _09791_ keymem.prev_key1_reg\[98\] _09790_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_110_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23519_ VGND VPWR VPWR VGND clk _00020_ reset_n keymem.key_mem\[14\]\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_135_363 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24499_ VGND VPWR VPWR VGND clk _00992_ reset_n keymem.key_mem\[9\]\[108\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_11_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17040_ VGND VPWR VPWR VGND _03084_ keymem.key_mem\[14\]\[61\] _03162_ _03163_ sky130_fd_sc_hd__mux2_2
XFILLER_0_145_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14252_ VGND VPWR VPWR VGND _09718_ _09716_ _09723_ _09722_ _09720_ sky130_fd_sc_hd__o211a_2
XFILLER_0_40_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_21_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_85_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13203_ VGND VPWR VGND VPWR _08016_ keymem.key_mem\[7\]\[103\] _08700_ _08702_ _08703_
+ _07573_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_180_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14183_ VGND VPWR VGND VPWR _09654_ _09651_ _09105_ _09652_ _09653_ sky130_fd_sc_hd__a211o_2
XFILLER_0_81_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_556 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_46_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13134_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[96\] _08124_ _08640_ _08636_ _08641_
+ sky130_fd_sc_hd__o22a_2
X_18991_ VGND VPWR _04822_ enc_block.block_w3_reg\[17\] enc_block.block_w1_reg\[1\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_81_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17942_ VGND VPWR _00245_ _03892_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13065_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[90\] _07652_ keymem.key_mem\[8\]\[90\]
+ _08211_ _08578_ sky130_fd_sc_hd__a22o_2
XFILLER_0_29_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1032 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_256_1309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12016_ VGND VPWR _07618_ _07602_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_178_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17873_ VGND VPWR _00223_ _03845_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_206_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_121_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19612_ VGND VPWR VPWR VGND _05205_ _05031_ keymem.key_mem\[12\]\[99\] _05209_ sky130_fd_sc_hd__mux2_2
X_16824_ VGND VPWR VPWR VGND _10820_ _10821_ _02864_ _02966_ sky130_fd_sc_hd__or3_2
XFILLER_0_254_1022 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_92_2_Right_164 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_254_1033 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_156_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_205_356 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19543_ VGND VPWR _00566_ _05172_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_92_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16755_ VGND VPWR _02904_ _02903_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_152_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13967_ VGND VPWR VPWR VGND _09298_ _09266_ _09296_ _09439_ sky130_fd_sc_hd__or3_2
XFILLER_0_156_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15706_ enc_block.sword_ctr_reg\[1\] _11162_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[18\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_92_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19474_ VPWR VGND keymem.key_mem\[12\]\[34\] _05136_ _05128_ VPWR VGND sky130_fd_sc_hd__and2_2
X_12918_ VPWR VGND VPWR VGND _08445_ keymem.key_mem\[12\]\[75\] _07722_ keymem.key_mem\[8\]\[75\]
+ _08265_ _08446_ sky130_fd_sc_hd__a221o_2
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16686_ VGND VPWR VPWR VGND _02662_ keymem.key_mem\[14\]\[30\] _02839_ _02840_ sky130_fd_sc_hd__mux2_2
X_13898_ VPWR VGND VGND VPWR _09331_ _09370_ _09319_ sky130_fd_sc_hd__nor2_2
XFILLER_0_5_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18425_ VPWR VGND VGND VPWR _04313_ enc_block.round_key\[64\] _04311_ sky130_fd_sc_hd__nand2_2
XFILLER_0_9_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15637_ VGND VPWR _09721_ key[14] _11095_ _09719_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_12849_ VGND VPWR VGND VPWR _08384_ _07712_ keymem.key_mem\[6\]\[68\] _08381_ _08383_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_232_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18356_ VPWR VGND VGND VPWR _04252_ _03996_ _04250_ sky130_fd_sc_hd__nand2_2
XFILLER_0_229_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15568_ VGND VPWR VGND VPWR _11025_ _11024_ _11027_ _11026_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_90_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17307_ VGND VPWR _00100_ _03402_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14519_ VGND VPWR _09988_ _09987_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18287_ VGND VPWR _04190_ _03973_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_4_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15499_ VPWR VGND VGND VPWR _10648_ _10706_ _10957_ _10958_ _10959_ sky130_fd_sc_hd__and4b_2
XFILLER_0_43_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17238_ VGND VPWR _00093_ _03340_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_163_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_821 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_163_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17169_ VGND VPWR _03279_ _03278_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_261_1059 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_180 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_243_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20180_ VGND VPWR _00865_ _05510_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_86_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_12_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_898 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_229_949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_204_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_161_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_228_448 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_196_1201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_237_960 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_100_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_193_21 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23870_ VGND VPWR VPWR VGND clk _00363_ reset_n enc_block.block_w2_reg\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_98_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_100_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22821_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[120\] _06860_ _06859_ _05075_ _02156_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_135_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_170_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25540_ VGND VPWR VPWR VGND clk _02033_ reset_n keymem.key_mem\[1\]\[125\] sky130_fd_sc_hd__dfrtp_2
X_22752_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[70\] _06837_ _06836_ _04983_ _02106_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_17_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21703_ VGND VPWR VPWR VGND _06319_ _03090_ keymem.key_mem\[4\]\[54\] _06321_ sky130_fd_sc_hd__mux2_2
X_25471_ VGND VPWR VPWR VGND clk _01964_ reset_n keymem.key_mem\[1\]\[56\] sky130_fd_sc_hd__dfrtp_2
X_22683_ VGND VPWR _02065_ _06813_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_250_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24422_ VGND VPWR VPWR VGND clk _00915_ reset_n keymem.key_mem\[9\]\[31\] sky130_fd_sc_hd__dfrtp_2
X_21634_ VGND VPWR _01545_ _06284_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_111_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24353_ VGND VPWR VPWR VGND clk _00846_ reset_n keymem.key_mem\[10\]\[90\] sky130_fd_sc_hd__dfrtp_2
X_21565_ VGND VPWR VPWR VGND _06242_ _03607_ keymem.key_mem\[5\]\[118\] _06247_ sky130_fd_sc_hd__mux2_2
XFILLER_0_132_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_7_583 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23304_ VGND VPWR _07185_ enc_block.block_w0_reg\[18\] _07184_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20516_ VGND VPWR _01022_ _05689_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24284_ VGND VPWR VPWR VGND clk _00777_ reset_n keymem.key_mem\[10\]\[21\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_181_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21496_ VGND VPWR VPWR VGND _06209_ _03374_ keymem.key_mem\[5\]\[85\] _06211_ sky130_fd_sc_hd__mux2_2
XFILLER_0_132_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_372 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23235_ _07121_ _07123_ _04103_ _07122_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_181_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1130 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20447_ VGND VPWR _00990_ _05652_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_30_320 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23166_ VGND VPWR VPWR VGND _07054_ _03599_ keymem.prev_key1_reg\[117\] _07068_ sky130_fd_sc_hd__mux2_2
XFILLER_0_222_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20378_ VGND VPWR _00957_ _05616_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_247_735 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22117_ VGND VPWR VPWR VGND _06538_ _05073_ keymem.key_mem\[3\]\[119\] _06542_ sky130_fd_sc_hd__mux2_2
XFILLER_0_63_1098 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_222_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23097_ VGND VPWR VPWR VGND _06992_ _07024_ keymem.prev_key1_reg\[91\] _07025_ sky130_fd_sc_hd__mux2_2
X_22048_ VGND VPWR VPWR VGND _06494_ _05010_ keymem.key_mem\[3\]\[86\] _06506_ sky130_fd_sc_hd__mux2_2
XFILLER_0_206_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_238_1028 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_237_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14870_ VGND VPWR VGND VPWR _10334_ _10221_ _10335_ _09821_ _09703_ sky130_fd_sc_hd__nand4_2
X_13821_ VGND VPWR _09293_ _09292_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25807_ keymem.prev_key1_reg\[123\] clk _02300_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_203_827 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_255_1386 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1228 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23999_ VGND VPWR VPWR VGND clk _00492_ reset_n keymem.key_mem\[13\]\[120\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_15_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16540_ _09589_ _02699_ keymem.round_ctr_reg\[0\] _09629_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_138_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13752_ VPWR VGND VGND VPWR _09221_ _09222_ _09224_ _09223_ _09080_ sky130_fd_sc_hd__o22ai_2
X_25738_ keymem.prev_key1_reg\[54\] clk _02231_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_253_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12703_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[54\] _07716_ keymem.key_mem\[12\]\[54\]
+ _07620_ _08252_ sky130_fd_sc_hd__a22o_2
X_16471_ VGND VPWR VGND VPWR _11249_ _11257_ _11313_ _11307_ _02632_ sky130_fd_sc_hd__o22a_2
X_13683_ VGND VPWR VGND VPWR _09153_ _09122_ _09154_ _09132_ _09155_ sky130_fd_sc_hd__o22a_2
X_25669_ VGND VPWR VPWR VGND clk _02162_ reset_n keymem.key_mem\[0\]\[126\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_214_1083 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18210_ VGND VPWR _04119_ enc_block.block_w1_reg\[21\] _04118_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15422_ VGND VPWR VGND VPWR _10566_ _10751_ _10593_ _10618_ _10883_ sky130_fd_sc_hd__o22a_2
XFILLER_0_6_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12634_ VGND VPWR VGND VPWR _08190_ _08150_ keymem.key_mem\[3\]\[47\] _08187_ _08189_
+ sky130_fd_sc_hd__a211o_2
X_19190_ VGND VPWR VGND VPWR _04960_ keymem.key_mem_we _03083_ _04924_ _00425_ sky130_fd_sc_hd__a31o_2
XFILLER_0_31_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_18141_ VGND VPWR _04056_ _04054_ _04055_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_38_497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15353_ _10775_ _10815_ keymem.round_ctr_reg\[0\] _10814_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_0_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12565_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[41\] _07918_ keymem.key_mem\[11\]\[41\]
+ _07658_ _08127_ sky130_fd_sc_hd__a22o_2
X_14304_ VGND VPWR VGND VPWR _09466_ _09441_ _09559_ _09408_ _09774_ sky130_fd_sc_hd__o22a_2
XFILLER_0_53_456 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_108_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18072_ VGND VPWR _03993_ _03973_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_262_1313 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15284_ VGND VPWR _10747_ _10746_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_41_629 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12496_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[34\] _07893_ _08064_ _08060_ _08065_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_184_1171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_149_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17023_ VPWR VGND VPWR VGND _03147_ key[188] _10322_ sky130_fd_sc_hd__or2_2
X_14235_ VGND VPWR _09106_ _09704_ _09706_ _09705_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_150_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14166_ VGND VPWR _09637_ _07378_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_145_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13117_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[95\] _07872_ keymem.key_mem\[1\]\[95\]
+ _07624_ _08625_ sky130_fd_sc_hd__a22o_2
XFILLER_0_238_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18974_ VPWR VGND _04807_ enc_block.block_w0_reg\[14\] enc_block.block_w1_reg\[7\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_14097_ VPWR VGND VGND VPWR _09480_ _09352_ _09568_ _09327_ _09391_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_226_908 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_221_1076 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17925_ VGND VPWR VPWR VGND _03876_ key[227] keymem.prev_key1_reg\[99\] _03881_ sky130_fd_sc_hd__mux2_2
X_13048_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[88\] _07924_ keymem.key_mem\[4\]\[88\]
+ _08077_ _08563_ sky130_fd_sc_hd__a22o_2
XFILLER_0_253_749 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_193_1418 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_147_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17856_ VGND VPWR VPWR VGND _03814_ _03833_ keymem.prev_key0_reg\[77\] _03834_ sky130_fd_sc_hd__mux2_2
XFILLER_0_206_654 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16807_ VGND VPWR VPWR VGND _09521_ key[168] keymem.prev_key1_reg\[40\] _02951_ sky130_fd_sc_hd__mux2_2
XFILLER_0_156_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17787_ VGND VPWR VGND VPWR _03737_ keymem.prev_key1_reg\[56\] _03679_ _03786_ sky130_fd_sc_hd__a21o_2
X_14999_ VGND VPWR _10463_ _10452_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_93_2_Right_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_117_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16738_ VGND VPWR VPWR VGND _09793_ _02887_ _02886_ _02888_ sky130_fd_sc_hd__mux2_2
X_19526_ VGND VPWR VGND VPWR _05163_ keymem.key_mem_we _03130_ _05135_ _00558_ sky130_fd_sc_hd__a31o_2
XFILLER_0_163_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_156_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_729 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_53_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19457_ VGND VPWR VGND VPWR _05126_ keymem.key_mem_we _02743_ _05121_ _00526_ sky130_fd_sc_hd__a31o_2
XFILLER_0_5_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16669_ VPWR VGND VGND VPWR _02823_ _02817_ _02822_ sky130_fd_sc_hd__nand2_2
XFILLER_0_8_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_902 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18408_ VPWR VGND VPWR VGND _04298_ block[127] _04213_ enc_block.block_w0_reg\[31\]
+ _04276_ _04299_ sky130_fd_sc_hd__a221o_2
XFILLER_0_5_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19388_ VGND VPWR _00497_ _05086_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_88_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_401 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18339_ _04235_ _04237_ _04008_ _04236_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_267_1257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21350_ VGND VPWR _01411_ _06134_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_71_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_163_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20301_ VGND VPWR VPWR VGND _05569_ _02924_ keymem.key_mem\[9\]\[37\] _05576_ sky130_fd_sc_hd__mux2_2
XFILLER_0_167_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21281_ VGND VPWR _01380_ _06096_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_163_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_640 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_128_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23020_ VGND VPWR _02236_ _06979_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_4_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20232_ VGND VPWR VPWR VGND _05535_ _10099_ keymem.key_mem\[9\]\[4\] _05540_ sky130_fd_sc_hd__mux2_2
XFILLER_0_124_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20163_ VGND VPWR _00857_ _05501_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_25_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_216_407 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_99_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20094_ VGND VPWR _05465_ _03227_ _00824_ _05402_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_24971_ VGND VPWR VPWR VGND clk _01464_ reset_n keymem.key_mem\[5\]\[68\] sky130_fd_sc_hd__dfrtp_2
X_23922_ VGND VPWR VPWR VGND clk _00415_ reset_n keymem.key_mem\[13\]\[43\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23853_ VGND VPWR VPWR VGND clk _00346_ reset_n enc_block.block_w2_reg\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_174_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_212_624 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_79_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_135_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22804_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[105\] _06858_ _06857_ _05043_ _02141_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_174_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23784_ VGND VPWR VPWR VGND clk _00277_ reset_n enc_block.block_w0_reg\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_71_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_977 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20996_ VGND VPWR VPWR VGND _05945_ _05045_ keymem.key_mem\[7\]\[106\] _05946_ sky130_fd_sc_hd__mux2_2
XFILLER_0_135_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25523_ VGND VPWR VPWR VGND clk _02016_ reset_n keymem.key_mem\[1\]\[108\] sky130_fd_sc_hd__dfrtp_2
X_22735_ VGND VPWR _02098_ _06832_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_71_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25454_ VGND VPWR VPWR VGND clk _01947_ reset_n keymem.key_mem\[1\]\[39\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_109_138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22666_ VGND VPWR _02057_ _06804_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_164_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_935 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24405_ VGND VPWR VPWR VGND clk _00898_ reset_n keymem.key_mem\[9\]\[14\] sky130_fd_sc_hd__dfrtp_2
X_21617_ VGND VPWR VPWR VGND _06275_ _11039_ keymem.key_mem\[4\]\[13\] _06276_ sky130_fd_sc_hd__mux2_2
X_25385_ VGND VPWR VPWR VGND clk _01878_ reset_n keymem.key_mem\[2\]\[98\] sky130_fd_sc_hd__dfrtp_2
X_22597_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[109\] _06775_ _06774_ _05052_ _02017_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_8_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1075 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_62_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24336_ VGND VPWR VPWR VGND clk _00829_ reset_n keymem.key_mem\[10\]\[73\] sky130_fd_sc_hd__dfrtp_2
X_12350_ VPWR VGND VPWR VGND _07931_ keymem.key_mem\[11\]\[21\] _07600_ keymem.key_mem\[1\]\[21\]
+ _07799_ _07932_ sky130_fd_sc_hd__a221o_2
XFILLER_0_51_927 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21548_ VGND VPWR VPWR VGND _06231_ _03555_ keymem.key_mem\[5\]\[110\] _06238_ sky130_fd_sc_hd__mux2_2
XFILLER_0_23_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_1496 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_990 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12281_ VPWR VGND VPWR VGND _07867_ keymem.key_mem\[13\]\[16\] _07587_ keymem.key_mem\[3\]\[16\]
+ _07618_ _07868_ sky130_fd_sc_hd__a221o_2
XFILLER_0_107_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21479_ VGND VPWR VPWR VGND _06196_ _03306_ keymem.key_mem\[5\]\[77\] _06202_ sky130_fd_sc_hd__mux2_2
X_24267_ VGND VPWR VPWR VGND clk _00760_ reset_n keymem.key_mem\[10\]\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_146_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14020_ VGND VPWR VGND VPWR _09491_ _09490_ _09492_ _09488_ _09484_ sky130_fd_sc_hd__nand4_2
XFILLER_0_31_651 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23218_ VPWR VGND _07107_ enc_block.block_w1_reg\[10\] enc_block.block_w2_reg\[1\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_31_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24198_ VGND VPWR VPWR VGND clk _00691_ reset_n keymem.key_mem\[11\]\[63\] sky130_fd_sc_hd__dfrtp_2
X_23149_ VGND VPWR _02286_ _07058_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_219_234 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_43_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15971_ _11174_ _11427_ _11233_ _11247_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_179_1251 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_257_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17710_ VGND VPWR VPWR VGND _03729_ _03739_ _02717_ _03740_ sky130_fd_sc_hd__or3_2
XFILLER_0_41_1193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14922_ VGND VPWR _10386_ _09717_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18690_ VPWR VGND VPWR VGND _04551_ _04550_ _04549_ enc_block.block_w1_reg\[26\]
+ _04328_ _00334_ sky130_fd_sc_hd__a221o_2
XFILLER_0_26_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17641_ VGND VPWR VPWR VGND _03681_ _03689_ keymem.prev_key0_reg\[6\] _03690_ sky130_fd_sc_hd__mux2_2
XFILLER_0_216_1101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_192_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14853_ VPWR VGND _10318_ _10317_ keymem.prev_key1_reg\[71\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_157_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13804_ enc_block.sword_ctr_reg\[1\] _09276_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[30\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_118_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_153_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17572_ VGND VPWR VPWR VGND _03593_ keymem.key_mem\[14\]\[122\] _03633_ _03634_ sky130_fd_sc_hd__mux2_2
X_14784_ VPWR VGND VPWR VGND _10067_ _10249_ _10121_ _09625_ _10250_ sky130_fd_sc_hd__or4_2
XFILLER_0_251_1058 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11996_ VGND VPWR _07599_ _07598_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_114_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19311_ VGND VPWR _00472_ _05034_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_15_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16523_ VPWR VGND _02683_ keymem.prev_key1_reg\[56\] keymem.prev_key1_reg\[24\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_153_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13735_ VPWR VGND VGND VPWR _09134_ _09207_ _09178_ sky130_fd_sc_hd__nor2_2
XFILLER_0_133_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_740 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_2_Left_582 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_85_356 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19242_ VPWR VGND VGND VPWR _04991_ keymem.key_mem\[13\]\[75\] _04880_ sky130_fd_sc_hd__nand2_2
X_16454_ VGND VPWR VGND VPWR _11282_ _11245_ _02615_ _11210_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_151_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13666_ VGND VPWR _09138_ _09137_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_6_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15405_ VGND VPWR VGND VPWR _10866_ _10562_ _10627_ _10543_ sky130_fd_sc_hd__o21a_2
X_12617_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[46\] _08050_ keymem.key_mem\[4\]\[46\]
+ _07665_ _08174_ sky130_fd_sc_hd__a22o_2
X_19173_ VGND VPWR VGND VPWR _04949_ keymem.key_mem_we _03025_ _04924_ _00419_ sky130_fd_sc_hd__a31o_2
XFILLER_0_5_306 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16385_ VGND VPWR VPWR VGND _02546_ _02545_ _02548_ _09722_ _02547_ sky130_fd_sc_hd__o211a_2
X_13597_ VGND VPWR _09069_ _09068_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_27_979 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18124_ VGND VPWR _04041_ _03973_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15336_ VGND VPWR VGND VPWR _10455_ _10797_ _10667_ _10583_ _10798_ sky130_fd_sc_hd__o22a_2
X_12548_ VPWR VGND VPWR VGND _08111_ keymem.key_mem\[13\]\[39\] _07730_ keymem.key_mem\[14\]\[39\]
+ _07963_ _08112_ sky130_fd_sc_hd__a221o_2
XFILLER_0_170_236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18055_ VGND VPWR _03976_ _03974_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_123_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15267_ VGND VPWR VGND VPWR _10666_ _07387_ _10729_ _10730_ sky130_fd_sc_hd__a21o_2
XFILLER_0_125_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12479_ VGND VPWR VGND VPWR _07542_ keymem.key_mem\[8\]\[33\] _08046_ _08048_ _08049_
+ _07663_ sky130_fd_sc_hd__a2111o_2
XPHY_EDGE_ROW_162_1_Left_429 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_164_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_111_314 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17006_ VGND VPWR _00070_ _03131_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14218_ VGND VPWR VGND VPWR _09145_ _09080_ _09221_ _09102_ _09689_ sky130_fd_sc_hd__o22a_2
XFILLER_0_125_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15198_ VGND VPWR _10662_ _10661_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_61_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_111_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14149_ VPWR VGND VPWR VGND _09618_ _09619_ _09620_ _09616_ _09617_ sky130_fd_sc_hd__or4b_2
XFILLER_0_61_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18957_ VGND VPWR _04792_ enc_block.block_w0_reg\[12\] enc_block.block_w0_reg\[13\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_201_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17908_ VGND VPWR VGND VPWR _03736_ keymem.prev_key0_reg\[93\] _03869_ _00234_ sky130_fd_sc_hd__a21o_2
X_18888_ _04728_ _04730_ _04727_ _04729_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_17839_ VGND VPWR _00212_ _03822_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_174_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_410 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_178_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_233_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_955 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20850_ VPWR VGND keymem.key_mem\[7\]\[37\] _05869_ _05856_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_171_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_2_Right_166 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_132_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19509_ VGND VPWR _00550_ _05154_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_190_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_212_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20781_ VGND VPWR VGND VPWR _05831_ keymem.key_mem_we _10194_ _05821_ _01145_ sky130_fd_sc_hd__a31o_2
XFILLER_0_18_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22520_ VGND VPWR _01968_ _06747_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_212_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_76_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_267_1021 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_91_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22451_ VGND VPWR _01927_ _06719_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_8_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_267_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21402_ VGND VPWR _01436_ _06161_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_44_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22382_ VGND VPWR _01895_ _06682_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25170_ VGND VPWR VPWR VGND clk _01663_ reset_n keymem.key_mem\[3\]\[11\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_114_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21333_ VGND VPWR _01403_ _06125_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24121_ VGND VPWR VPWR VGND clk _00614_ reset_n keymem.key_mem\[12\]\[114\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_161_269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_44_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_60_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1227 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_4_394 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24052_ VGND VPWR VPWR VGND clk _00545_ reset_n keymem.key_mem\[12\]\[45\] sky130_fd_sc_hd__dfrtp_2
X_21264_ VGND VPWR VPWR VGND _06087_ _03518_ keymem.key_mem\[6\]\[104\] _06088_ sky130_fd_sc_hd__mux2_2
XFILLER_0_13_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_198_1104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23003_ VGND VPWR _02229_ _06969_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20215_ VGND VPWR _00882_ _05528_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_187_2_Left_658 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21195_ VGND VPWR _01339_ _06051_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_99_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20146_ VGND VPWR _00849_ _05492_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_204_1093 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_99_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_216_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_216_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24954_ VGND VPWR VPWR VGND clk _01447_ reset_n keymem.key_mem\[5\]\[51\] sky130_fd_sc_hd__dfrtp_2
X_20077_ VGND VPWR _00816_ _05456_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_235_1009 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23905_ VGND VPWR VPWR VGND clk _00398_ reset_n keymem.key_mem\[13\]\[26\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_197_612 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24885_ VGND VPWR VPWR VGND clk _01378_ reset_n keymem.key_mem\[6\]\[110\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_234_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11850_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[28\] dec_new_block\[92\]
+ _07489_ sky130_fd_sc_hd__mux2_2
X_23836_ VGND VPWR VPWR VGND clk _00329_ reset_n enc_block.block_w1_reg\[21\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_252_1367 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11781_ VGND VPWR result[57] _07454_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_94_120 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23767_ keymem.prev_key0_reg\[123\] clk _00264_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_36_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20979_ VGND VPWR VPWR VGND _05934_ _05029_ keymem.key_mem\[7\]\[98\] _05937_ sky130_fd_sc_hd__mux2_2
X_13520_ VPWR VGND VGND VPWR enc_block.block_w1_reg\[4\] enc_block.sword_ctr_reg\[0\]
+ _08992_ sky130_fd_sc_hd__or2b_2
XFILLER_0_71_1175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25506_ VGND VPWR VPWR VGND clk _01999_ reset_n keymem.key_mem\[1\]\[91\] sky130_fd_sc_hd__dfrtp_2
X_22718_ VGND VPWR _02089_ _06824_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_3_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23698_ keymem.prev_key0_reg\[54\] clk _00195_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_211_1086 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25437_ VGND VPWR VPWR VGND clk _01930_ reset_n keymem.key_mem\[1\]\[22\] sky130_fd_sc_hd__dfrtp_2
X_13451_ VGND VPWR VGND VPWR _07370_ result_valid _07368_ _00011_ sky130_fd_sc_hd__a21o_2
XFILLER_0_3_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22649_ VGND VPWR _02049_ _06795_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_152_214 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12402_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[26\] _07865_ keymem.key_mem\[12\]\[26\]
+ _07621_ _07979_ sky130_fd_sc_hd__a22o_2
X_16170_ VGND VPWR _11624_ _09516_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_1_1260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25368_ VGND VPWR VPWR VGND clk _01861_ reset_n keymem.key_mem\[2\]\[81\] sky130_fd_sc_hd__dfrtp_2
X_13382_ VPWR VGND VPWR VGND _08863_ keymem.key_mem\[6\]\[121\] _07711_ keymem.key_mem\[8\]\[121\]
+ _08265_ _08864_ sky130_fd_sc_hd__a221o_2
XFILLER_0_24_938 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_23_426 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15121_ VGND VPWR VGND VPWR _10585_ _10584_ _10515_ _10465_ sky130_fd_sc_hd__o21a_2
X_24319_ VGND VPWR VPWR VGND clk _00812_ reset_n keymem.key_mem\[10\]\[56\] sky130_fd_sc_hd__dfrtp_2
X_12333_ VPWR VGND VPWR VGND _07915_ keymem.key_mem\[11\]\[20\] _07912_ keymem.key_mem\[12\]\[20\]
+ _07808_ _07916_ sky130_fd_sc_hd__a221o_2
X_25299_ VGND VPWR VPWR VGND clk _01792_ reset_n keymem.key_mem\[2\]\[12\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_51_779 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_107_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15052_ VGND VPWR VGND VPWR _10516_ _10500_ _10514_ _10440_ _10477_ sky130_fd_sc_hd__a211o_2
XFILLER_0_146_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12264_ VGND VPWR VGND VPWR _07786_ keymem.key_mem\[10\]\[15\] _07849_ _07851_ _07852_
+ _07663_ sky130_fd_sc_hd__a2111o_2
X_14003_ VGND VPWR _09475_ _09474_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_43_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_852 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19860_ VGND VPWR VPWR VGND _05339_ keymem.key_mem\[11\]\[87\] _03393_ _05341_ sky130_fd_sc_hd__mux2_2
X_12195_ VGND VPWR _07788_ _07787_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_140_1_Right_741 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18811_ _04659_ _04661_ _04560_ _04660_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_207_204 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_78_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19791_ VGND VPWR VPWR VGND _05303_ keymem.key_mem\[11\]\[54\] _03091_ _05305_ sky130_fd_sc_hd__mux2_2
XFILLER_0_263_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15954_ VGND VPWR VGND VPWR _11410_ _11407_ _11287_ _11409_ _11408_ _11224_ sky130_fd_sc_hd__a32o_2
X_18742_ VPWR VGND _04598_ _04597_ enc_block.round_key\[32\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_37_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14905_ VGND VPWR VPWR VGND _09864_ keymem.key_mem\[14\]\[7\] _10369_ _10370_ sky130_fd_sc_hd__mux2_2
X_18673_ VGND VPWR _04536_ enc_block.block_w2_reg\[17\] _04469_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_15885_ _11339_ _11341_ _11338_ _11340_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_14836_ VPWR VGND VGND VPWR _09302_ _10301_ _09582_ sky130_fd_sc_hd__nor2_2
X_17624_ VGND VPWR VPWR VGND _03675_ _03677_ keymem.prev_key0_reg\[1\] _03678_ sky130_fd_sc_hd__mux2_2
XFILLER_0_118_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_114_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17555_ VPWR VGND VGND VPWR keylen _03617_ _03618_ _03619_ sky130_fd_sc_hd__nor3_2
XFILLER_0_15_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14767_ VGND VPWR VPWR VGND _10126_ _10232_ _09902_ _10233_ sky130_fd_sc_hd__or3_2
X_11979_ VGND VPWR _07582_ _07581_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_19_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16506_ VGND VPWR VGND VPWR _09505_ _09429_ _02666_ _10360_ sky130_fd_sc_hd__a21oi_2
X_13718_ VPWR VGND VGND VPWR _09010_ _09190_ _09057_ sky130_fd_sc_hd__nor2_2
XFILLER_0_89_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17486_ VPWR VGND _09533_ _03559_ _03558_ VPWR VGND sky130_fd_sc_hd__and2_2
X_14698_ VPWR VGND VGND VPWR _09103_ _09221_ _09114_ _09091_ _10165_ _10164_ sky130_fd_sc_hd__o221a_2
XFILLER_0_89_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16437_ VGND VPWR VGND VPWR _02598_ _02597_ _02599_ keymem.prev_key1_reg\[86\] sky130_fd_sc_hd__a21oi_2
X_19225_ VPWR VGND VGND VPWR _04981_ keymem.key_mem\[13\]\[68\] _04880_ sky130_fd_sc_hd__nand2_2
X_13649_ VGND VPWR _09121_ _09120_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_143_203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19156_ VGND VPWR _00413_ _04938_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16368_ VGND VPWR VGND VPWR _11372_ _11305_ _02531_ _11404_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_26_275 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_724 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18107_ VPWR VGND _04025_ _04024_ enc_block.block_w2_reg\[12\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15319_ VPWR VGND VGND VPWR _10587_ _10781_ _10414_ sky130_fd_sc_hd__nor2_2
XFILLER_0_87_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19087_ VPWR VGND keymem.key_mem\[13\]\[13\] _04898_ _04887_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16299_ VGND VPWR VGND VPWR _02461_ _02460_ _02462_ _02463_ sky130_fd_sc_hd__a21o_2
XFILLER_0_227_1060 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_42_779 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1019 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18038_ VPWR VGND _03960_ enc_block.block_w0_reg\[31\] enc_block.block_w0_reg\[24\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_125_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_876 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_65_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_375 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_199_1446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_22_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20000_ VGND VPWR _00779_ _05416_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_199_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_676 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19989_ VGND VPWR _00774_ _05410_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_94_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_1085 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21951_ VGND VPWR _01692_ _06454_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_55_1104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_222_741 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20902_ VGND VPWR VGND VPWR _05896_ keymem.key_mem_we _03162_ _05893_ _01201_ sky130_fd_sc_hd__a31o_2
X_24670_ VGND VPWR VPWR VGND clk _01163_ reset_n keymem.key_mem\[7\]\[23\] sky130_fd_sc_hd__dfrtp_2
X_21882_ VPWR VGND keymem.key_mem\[3\]\[9\] _06417_ _06413_ VPWR VGND sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_19_Left_287 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_136_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23621_ VGND VPWR VPWR VGND clk _00122_ reset_n keymem.key_mem\[14\]\[110\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_72_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20833_ VGND VPWR VGND VPWR _05859_ keymem.key_mem_we _02812_ _05850_ _01169_ sky130_fd_sc_hd__a31o_2
XFILLER_0_33_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_120 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_95_2_Right_167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_204_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_134_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23552_ VGND VPWR VPWR VGND clk _00053_ reset_n keymem.key_mem\[14\]\[41\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20764_ VGND VPWR _05820_ _05819_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22503_ VGND VPWR VPWR VGND _06739_ keymem.key_mem\[1\]\[51\] _03068_ _06740_ sky130_fd_sc_hd__mux2_2
XFILLER_0_193_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23483_ VGND VPWR _07345_ _07343_ _07344_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_20695_ VGND VPWR _05783_ _05675_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_247_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25222_ VGND VPWR VPWR VGND clk _01715_ reset_n keymem.key_mem\[3\]\[63\] sky130_fd_sc_hd__dfrtp_2
X_22434_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[11\] _06707_ _06706_ _04894_ _01919_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_91_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_91 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25153_ VGND VPWR VPWR VGND clk _01646_ reset_n keymem.key_mem\[4\]\[122\] sky130_fd_sc_hd__dfrtp_2
X_22365_ VGND VPWR _01887_ _06673_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_28_Left_296 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24104_ VGND VPWR VPWR VGND clk _00597_ reset_n keymem.key_mem\[12\]\[97\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_108_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21316_ VGND VPWR _06116_ _06115_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_143_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25084_ VGND VPWR VPWR VGND clk _01577_ reset_n keymem.key_mem\[4\]\[53\] sky130_fd_sc_hd__dfrtp_2
X_22296_ VGND VPWR _06637_ _03279_ _01854_ _06567_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_142_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21247_ VGND VPWR VPWR VGND _06076_ _03466_ keymem.key_mem\[6\]\[96\] _06079_ sky130_fd_sc_hd__mux2_2
X_24035_ VGND VPWR VPWR VGND clk _00528_ reset_n keymem.key_mem\[12\]\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_206_1199 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_264_619 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21178_ VGND VPWR VPWR VGND _06040_ _03183_ keymem.key_mem\[6\]\[63\] _06043_ sky130_fd_sc_hd__mux2_2
XFILLER_0_257_682 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_256_170 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_258_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20129_ VGND VPWR VPWR VGND _05482_ _03374_ keymem.key_mem\[10\]\[85\] _05484_ sky130_fd_sc_hd__mux2_2
XFILLER_0_245_866 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_219_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_258_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_719 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_254_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24937_ VGND VPWR VPWR VGND clk _01430_ reset_n keymem.key_mem\[5\]\[34\] sky130_fd_sc_hd__dfrtp_2
X_12951_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[78\] _08124_ _08475_ _08469_ _08476_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_260_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11902_ VGND VPWR VPWR VGND encdec enc_block.block_w0_reg\[22\] dec_new_block\[118\]
+ _07515_ sky130_fd_sc_hd__mux2_2
X_15670_ VGND VPWR VGND VPWR _10627_ _10538_ _10609_ _10530_ _11127_ sky130_fd_sc_hd__o22a_2
XFILLER_0_213_752 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_115_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24868_ VGND VPWR VPWR VGND clk _01361_ reset_n keymem.key_mem\[6\]\[93\] sky130_fd_sc_hd__dfrtp_2
X_12882_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[72\] _07588_ keymem.key_mem\[2\]\[72\]
+ _07816_ _08413_ sky130_fd_sc_hd__a22o_2
XFILLER_0_154_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14621_ VGND VPWR _10089_ keymem.prev_key1_reg\[68\] _10088_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_11833_ VGND VPWR result[83] _07480_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23819_ VGND VPWR VPWR VGND clk _00312_ reset_n enc_block.block_w1_reg\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_115_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24799_ VGND VPWR VPWR VGND clk _01292_ reset_n keymem.key_mem\[6\]\[24\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_114_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_197_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17340_ VPWR VGND VGND VPWR _11456_ _03432_ key[220] sky130_fd_sc_hd__nor2_2
X_14552_ VGND VPWR VGND VPWR _09188_ _09059_ _09179_ _10020_ sky130_fd_sc_hd__a21o_2
XFILLER_0_261_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11764_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[17\] dec_new_block\[49\]
+ _07446_ sky130_fd_sc_hd__mux2_2
X_13503_ VPWR VGND VPWR VGND _08974_ _08948_ _08973_ _08945_ enc_block.block_w2_reg\[7\]
+ _08975_ sky130_fd_sc_hd__a221o_2
X_17271_ VGND VPWR VGND VPWR _03370_ _03302_ _02927_ key[85] sky130_fd_sc_hd__o21a_2
X_14483_ VGND VPWR VGND VPWR _09221_ _09109_ _09090_ _09127_ _09952_ sky130_fd_sc_hd__o22a_2
XFILLER_0_55_348 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_82_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_165_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11695_ VGND VPWR result[14] _07411_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19010_ VGND VPWR _04839_ _04780_ _04838_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_265_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16222_ VPWR VGND VGND VPWR _11482_ _11466_ _02387_ _11420_ _11400_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_125_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13434_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[126\] _08027_ _08910_ _08906_ _08911_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_64_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_226_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_521 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16153_ VPWR VGND VGND VPWR _11607_ _11606_ _11605_ _11603_ _11345_ _11246_ sky130_fd_sc_hd__o2111a_2
X_13365_ VGND VPWR enc_block.round_key\[119\] _08848_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15104_ VGND VPWR VPWR VGND _10440_ _10466_ _10451_ _10568_ sky130_fd_sc_hd__or3_2
X_12316_ VPWR VGND VPWR VGND _07899_ keymem.key_mem\[5\]\[19\] _07779_ keymem.key_mem\[13\]\[19\]
+ _07622_ _07900_ sky130_fd_sc_hd__a221o_2
XFILLER_0_80_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16084_ VGND VPWR VGND VPWR _11536_ _11535_ _11537_ _11539_ sky130_fd_sc_hd__a21o_2
X_13296_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[113\] _07782_ keymem.key_mem\[10\]\[113\]
+ _07785_ _08786_ sky130_fd_sc_hd__a22o_2
XFILLER_0_32_790 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_122_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15035_ VPWR VGND VGND VPWR _10498_ _10499_ _10496_ sky130_fd_sc_hd__nor2_2
X_19912_ VGND VPWR VPWR VGND _05361_ keymem.key_mem\[11\]\[112\] _03567_ _05368_ sky130_fd_sc_hd__mux2_2
XFILLER_0_43_1030 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12247_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[14\] _07835_ keymem.key_mem\[1\]\[14\]
+ _07800_ _07836_ sky130_fd_sc_hd__a22o_2
XFILLER_0_20_974 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_141_1_Right_742 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19843_ VGND VPWR VPWR VGND _05328_ keymem.key_mem\[11\]\[79\] _03322_ _05332_ sky130_fd_sc_hd__mux2_2
XFILLER_0_236_822 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12178_ VPWR VGND VPWR VGND keymem.key_mem\[4\]\[9\] _07636_ keymem.key_mem\[1\]\[9\]
+ _07624_ _07772_ sky130_fd_sc_hd__a22o_2
XFILLER_0_48_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19774_ VGND VPWR VPWR VGND _05292_ keymem.key_mem\[11\]\[46\] _03015_ _05296_ sky130_fd_sc_hd__mux2_2
XFILLER_0_236_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16986_ VGND VPWR VPWR VGND _03111_ _02691_ _03113_ _09514_ _03112_ sky130_fd_sc_hd__o211a_2
X_18725_ VPWR VGND VGND VPWR _04512_ _04583_ _04292_ sky130_fd_sc_hd__nor2_2
X_15937_ VPWR VGND VGND VPWR _11303_ _11320_ _11393_ _11352_ _11367_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_218_1037 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_194_1376 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_155_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15868_ VGND VPWR VPWR VGND _11265_ _11179_ _11233_ _11324_ sky130_fd_sc_hd__or3_2
X_18656_ VPWR VGND VPWR VGND _04521_ _04459_ _04520_ enc_block.block_w1_reg\[22\]
+ _04424_ _00330_ sky130_fd_sc_hd__a221o_2
XFILLER_0_259_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_118_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14819_ VGND VPWR VPWR VGND _09864_ keymem.key_mem\[14\]\[6\] _10284_ _10285_ sky130_fd_sc_hd__mux2_2
X_17607_ VGND VPWR VGND VPWR _03664_ _03302_ _08937_ key[127] sky130_fd_sc_hd__o21a_2
X_15799_ VPWR VGND VPWR VGND _11242_ _11254_ _11255_ _11220_ _11231_ sky130_fd_sc_hd__or4b_2
X_18587_ VPWR VGND VGND VPWR _04380_ _04460_ _04137_ sky130_fd_sc_hd__nor2_2
XFILLER_0_175_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_58_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17538_ VPWR VGND key[246] _03604_ _09523_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_171_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_89_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17469_ VGND VPWR _00120_ _03544_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_190_106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_412 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_89_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_1_Left_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19208_ VPWR VGND keymem.key_mem\[13\]\[61\] _04971_ _04961_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_13_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20480_ VGND VPWR _01006_ _05669_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_6_467 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_15_735 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_6_489 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_54_392 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19139_ VPWR VGND keymem.key_mem_we _04927_ _02913_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_242_1311 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_89_86 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22150_ VGND VPWR _01785_ _06560_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_278 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_749 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21101_ VGND VPWR _01294_ _06002_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_66_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22081_ VGND VPWR VPWR VGND _06516_ _05037_ keymem.key_mem\[3\]\[102\] _06523_ sky130_fd_sc_hd__mux2_2
XFILLER_0_1_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21032_ VGND VPWR _01263_ _05964_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_199_1254 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25840_ VGND VPWR VPWR VGND clk _02333_ reset_n enc_block.block_w3_reg\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_226_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_199_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25771_ keymem.prev_key1_reg\[87\] clk _02264_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22983_ VGND VPWR _02221_ _06957_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_242_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_198_239 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24722_ VGND VPWR VPWR VGND clk _01215_ reset_n keymem.key_mem\[7\]\[75\] sky130_fd_sc_hd__dfrtp_2
X_21934_ VGND VPWR VPWR VGND _06403_ _04922_ keymem.key_mem\[3\]\[33\] _06445_ sky130_fd_sc_hd__mux2_2
XFILLER_0_215_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24653_ VGND VPWR VPWR VGND clk _01146_ reset_n keymem.key_mem\[7\]\[6\] sky130_fd_sc_hd__dfrtp_2
X_21865_ VPWR VGND keymem.key_mem\[3\]\[1\] _06408_ _06406_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_49_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23604_ VGND VPWR VPWR VGND clk _00105_ reset_n keymem.key_mem\[14\]\[93\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_96_2_Right_168 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_132_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20816_ VGND VPWR _05850_ _05820_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24584_ VGND VPWR VPWR VGND clk _01077_ reset_n keymem.key_mem\[8\]\[65\] sky130_fd_sc_hd__dfrtp_2
X_21796_ VGND VPWR _01622_ _06369_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_37_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23535_ VGND VPWR VPWR VGND clk _00036_ reset_n keymem.key_mem\[14\]\[24\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_231_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20747_ VGND VPWR _01132_ _05810_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_247_1233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23466_ VPWR VGND VPWR VGND _07330_ _07117_ _07328_ sky130_fd_sc_hd__or2_2
XFILLER_0_68_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1244 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_36_Left_304 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_52_329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20678_ VGND VPWR _01099_ _05774_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_110_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25205_ VGND VPWR VPWR VGND clk _01698_ reset_n keymem.key_mem\[3\]\[46\] sky130_fd_sc_hd__dfrtp_2
X_22417_ VGND VPWR _06701_ _06695_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23397_ VPWR VGND VGND VPWR _07269_ _07265_ _07267_ sky130_fd_sc_hd__nand2_2
XFILLER_0_122_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13150_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[98\] _08090_ keymem.key_mem\[1\]\[98\]
+ _07558_ _08655_ sky130_fd_sc_hd__a22o_2
X_25136_ VGND VPWR VPWR VGND clk _01629_ reset_n keymem.key_mem\[4\]\[105\] sky130_fd_sc_hd__dfrtp_2
X_22348_ VGND VPWR _01879_ _06664_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_108_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12101_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[5\] _07631_ keymem.key_mem\[8\]\[5\]
+ _07654_ _07699_ sky130_fd_sc_hd__a22o_2
X_13081_ VPWR VGND VPWR VGND _08592_ keymem.key_mem\[3\]\[91\] _08009_ keymem.key_mem\[11\]\[91\]
+ _07902_ _08593_ sky130_fd_sc_hd__a221o_2
XFILLER_0_260_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_221_1428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25067_ VGND VPWR VPWR VGND clk _01560_ reset_n keymem.key_mem\[4\]\[36\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_108_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22279_ VGND VPWR _01846_ _06628_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_218_822 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24018_ VGND VPWR VPWR VGND clk _00511_ reset_n keymem.key_mem\[12\]\[11\] sky130_fd_sc_hd__dfrtp_2
X_12032_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[2\] _07586_ keymem.key_mem\[8\]\[2\]
+ _07539_ _07633_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_120_2_Left_591 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_217_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_79_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16840_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[75\] keymem.prev_key1_reg\[43\]
+ _02981_ _02980_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_45_Left_313 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_258_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_899 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_79_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16771_ VPWR VGND VGND VPWR _02918_ key[165] _09544_ sky130_fd_sc_hd__nand2_2
X_13983_ VPWR VGND VPWR VGND _09455_ _09446_ _09454_ sky130_fd_sc_hd__or2_2
XFILLER_0_191_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15722_ VPWR VGND VPWR VGND _11178_ enc_block.block_w0_reg\[17\] _09273_ sky130_fd_sc_hd__or2_2
X_18510_ VGND VPWR VGND VPWR _04389_ _04390_ _04316_ _04391_ enc_block.block_w1_reg\[7\]
+ sky130_fd_sc_hd__o2bb2a_2
X_12934_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[77\] _07724_ keymem.key_mem\[8\]\[77\]
+ _07540_ _08460_ sky130_fd_sc_hd__a22o_2
XFILLER_0_220_508 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_87_204 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19490_ VGND VPWR _00541_ _05144_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_16_Right_16 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18441_ VGND VPWR _04328_ _04314_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15653_ VPWR VGND _11110_ keymem.prev_key0_reg\[79\] keymem.prev_key0_reg\[47\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_119_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12865_ VPWR VGND VPWR VGND _08397_ keymem.key_mem\[14\]\[70\] _08003_ keymem.key_mem\[11\]\[70\]
+ _07781_ _08398_ sky130_fd_sc_hd__a221o_2
XPHY_EDGE_ROW_171_1_Left_438 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14604_ VGND VPWR VGND VPWR _10072_ _09574_ _09447_ _09876_ _10071_ sky130_fd_sc_hd__a211o_2
XFILLER_0_200_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11816_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[11\] dec_new_block\[75\]
+ _07472_ sky130_fd_sc_hd__mux2_2
X_18372_ VGND VPWR VGND VPWR _04265_ _04266_ _03974_ _04267_ enc_block.block_w0_reg\[27\]
+ sky130_fd_sc_hd__o2bb2a_2
X_15584_ VGND VPWR _00025_ _11042_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_189_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12796_ VGND VPWR VGND VPWR _07912_ keymem.key_mem\[11\]\[63\] _08333_ _08335_ _08336_
+ _08020_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_28_326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_95_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17323_ VPWR VGND VPWR VGND _03416_ _03413_ _03411_ key[218] _02723_ _03417_ sky130_fd_sc_hd__a221o_2
XFILLER_0_157_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14535_ VGND VPWR VPWR VGND _09996_ _10002_ _09119_ _10003_ sky130_fd_sc_hd__or3_2
XFILLER_0_141_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11747_ VGND VPWR result[40] _07437_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_44_808 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_54_Left_322 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_141_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_138_383 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17254_ VGND VPWR VGND VPWR _11151_ key[211] _03354_ _03355_ sky130_fd_sc_hd__a21o_2
X_14466_ VPWR VGND VGND VPWR _09099_ _09935_ _09036_ sky130_fd_sc_hd__nor2_2
XFILLER_0_4_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11678_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[6\] dec_new_block\[6\]
+ _07403_ sky130_fd_sc_hd__mux2_2
XFILLER_0_187_1180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16205_ VGND VPWR VPWR VGND _11345_ _11241_ _02370_ _02369_ _11387_ sky130_fd_sc_hd__o211a_2
XFILLER_0_226_1317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13417_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[125\] _07586_ keymem.key_mem\[3\]\[125\]
+ _07602_ _08895_ sky130_fd_sc_hd__a22o_2
XFILLER_0_10_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_543 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17185_ VGND VPWR VPWR VGND _03292_ _03293_ keymem.prev_key0_reg\[76\] _10327_ _10963_
+ sky130_fd_sc_hd__a31oi_2
XPHY_EDGE_ROW_25_Right_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14397_ VGND VPWR _09866_ _09523_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16136_ VPWR VGND VGND VPWR _11211_ _11590_ _11250_ sky130_fd_sc_hd__nor2_2
X_13348_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[118\] _07845_ keymem.key_mem\[1\]\[118\]
+ _07671_ _08833_ sky130_fd_sc_hd__a22o_2
XFILLER_0_267_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16067_ VPWR VGND VGND VPWR _11311_ _11522_ _11205_ sky130_fd_sc_hd__nor2_2
XFILLER_0_228_608 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_11_259 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13279_ VPWR VGND VPWR VGND _08770_ keymem.key_mem\[13\]\[111\] _07834_ keymem.key_mem\[8\]\[111\]
+ _07655_ _08771_ sky130_fd_sc_hd__a221o_2
XFILLER_0_23_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_227_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15018_ VGND VPWR _10482_ _10481_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_267_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1416 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_248_490 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_142_1_Right_743 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_97_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19826_ VGND VPWR VPWR VGND _05314_ keymem.key_mem\[11\]\[71\] _03252_ _05323_ sky130_fd_sc_hd__mux2_2
XFILLER_0_202_1394 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_237_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19757_ VGND VPWR VPWR VGND _05281_ keymem.key_mem\[11\]\[38\] _02934_ _05287_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_34_Right_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16969_ VPWR VGND VPWR VGND _03098_ _03095_ _02654_ _02655_ _03097_ _02496_ sky130_fd_sc_hd__o311a_2
XFILLER_0_237_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18708_ VPWR VGND VGND VPWR _04512_ _04568_ _04274_ sky130_fd_sc_hd__nor2_2
XFILLER_0_251_666 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_223_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_155_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19688_ VGND VPWR VPWR VGND _05247_ keymem.key_mem\[11\]\[5\] _10194_ _05251_ sky130_fd_sc_hd__mux2_2
XFILLER_0_91_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18639_ VPWR VGND _04506_ enc_block.block_w3_reg\[13\] enc_block.block_w3_reg\[12\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_148_114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_59_473 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_91_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21650_ VGND VPWR VPWR VGND _06286_ _02811_ keymem.key_mem\[4\]\[29\] _06293_ sky130_fd_sc_hd__mux2_2
XFILLER_0_8_1085 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_46_112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_136_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20601_ VGND VPWR VPWR VGND _05725_ _03067_ keymem.key_mem\[8\]\[51\] _05734_ sky130_fd_sc_hd__mux2_2
XFILLER_0_168_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21581_ VGND VPWR VPWR VGND _06116_ _03661_ keymem.key_mem\[5\]\[126\] _06255_ sky130_fd_sc_hd__mux2_2
XFILLER_0_7_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23320_ VPWR VGND VPWR VGND _07199_ block[11] _04139_ enc_block.block_w1_reg\[11\]
+ _03953_ _07200_ sky130_fd_sc_hd__a221o_2
X_20532_ VGND VPWR VPWR VGND _05692_ _02339_ keymem.key_mem\[8\]\[18\] _05698_ sky130_fd_sc_hd__mux2_2
XFILLER_0_144_331 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1220 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_28_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_144_353 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_6_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_776 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_244_1417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23251_ VGND VPWR VGND VPWR _07137_ _03949_ _04030_ _07138_ sky130_fd_sc_hd__a21o_2
XFILLER_0_209_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20463_ VGND VPWR VPWR VGND _05660_ _03580_ keymem.key_mem\[9\]\[114\] _05661_ sky130_fd_sc_hd__mux2_2
XFILLER_0_166_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22202_ VGND VPWR VPWR VGND _06578_ _02838_ keymem.key_mem\[2\]\[30\] _06588_ sky130_fd_sc_hd__mux2_2
XFILLER_0_63_1214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_63_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20394_ VGND VPWR _00965_ _05624_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23182_ VGND VPWR VPWR VGND _06880_ _07077_ keymem.prev_key1_reg\[123\] _07078_ sky130_fd_sc_hd__mux2_2
X_22133_ VGND VPWR VPWR VGND _06402_ _05089_ keymem.key_mem\[3\]\[127\] _06550_ sky130_fd_sc_hd__mux2_2
XFILLER_0_63_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_939 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22064_ VGND VPWR VPWR VGND _06494_ _05021_ keymem.key_mem\[3\]\[94\] _06514_ sky130_fd_sc_hd__mux2_2
XFILLER_0_10_270 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_206_Left_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21015_ VGND VPWR _01255_ _05955_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_52_Right_52 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_255_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25823_ VGND VPWR VPWR VGND clk _02316_ reset_n enc_block.block_w3_reg\[11\] sky130_fd_sc_hd__dfrtp_2
X_25754_ keymem.prev_key1_reg\[70\] clk _02247_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_202_508 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22966_ VGND VPWR _02214_ _06947_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_230_828 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_69_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24705_ VGND VPWR VPWR VGND clk _01198_ reset_n keymem.key_mem\[7\]\[58\] sky130_fd_sc_hd__dfrtp_2
X_21917_ VPWR VGND keymem.key_mem\[3\]\[25\] _06436_ _06427_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_179_261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25685_ keymem.prev_key1_reg\[1\] clk _02178_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_70_1218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_74_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22897_ VGND VPWR VPWR VGND _06878_ _10975_ keymem.prev_key1_reg\[12\] _06904_ sky130_fd_sc_hd__mux2_2
XFILLER_0_242_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12650_ VPWR VGND VPWR VGND _08203_ keymem.key_mem\[3\]\[49\] _07844_ keymem.key_mem\[8\]\[49\]
+ _07655_ _08204_ sky130_fd_sc_hd__a221o_2
X_24636_ VGND VPWR VPWR VGND clk _01129_ reset_n keymem.key_mem\[8\]\[117\] sky130_fd_sc_hd__dfrtp_2
X_21848_ VGND VPWR _01647_ _06396_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_77_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_210_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_139_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_215_Left_482 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_97_2_Right_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_808 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24567_ VGND VPWR VPWR VGND clk _01060_ reset_n keymem.key_mem\[8\]\[48\] sky130_fd_sc_hd__dfrtp_2
X_12581_ VPWR VGND VPWR VGND _08141_ keymem.key_mem\[14\]\[42\] _07963_ keymem.key_mem\[1\]\[42\]
+ _07901_ _08142_ sky130_fd_sc_hd__a221o_2
XFILLER_0_154_117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21779_ VGND VPWR _01614_ _06360_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_61_Right_61 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14320_ VPWR VGND VGND VPWR _09790_ _09759_ _09789_ sky130_fd_sc_hd__nand2_2
X_23518_ VGND VPWR VPWR VGND clk _00019_ reset_n keymem.key_mem\[14\]\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_53_638 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_110_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24498_ VGND VPWR VPWR VGND clk _00991_ reset_n keymem.key_mem\[9\]\[107\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_52_126 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_208_1003 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14251_ VGND VPWR _09722_ _09721_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_1369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23449_ VPWR VGND VPWR VGND _07314_ block[25] _03958_ enc_block.block_w3_reg\[25\]
+ _04504_ _07315_ sky130_fd_sc_hd__a221o_2
XFILLER_0_11_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13202_ VPWR VGND VPWR VGND _08701_ keymem.key_mem\[11\]\[103\] _07600_ keymem.key_mem\[1\]\[103\]
+ _07799_ _08702_ sky130_fd_sc_hd__a221o_2
XFILLER_0_81_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14182_ VGND VPWR VGND VPWR _09097_ _09094_ _09653_ _09156_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_145_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_81_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25119_ VGND VPWR VPWR VGND clk _01612_ reset_n keymem.key_mem\[4\]\[88\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_238_906 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13133_ VGND VPWR VGND VPWR _08640_ _07968_ keymem.key_mem\[9\]\[96\] _08637_ _08639_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_42_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_103_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18990_ VPWR VGND VPWR VGND _04821_ _04788_ _04820_ enc_block.block_w2_reg\[24\]
+ _04613_ _00364_ sky130_fd_sc_hd__a221o_2
XFILLER_0_29_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_224_Left_491 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17941_ VGND VPWR VPWR VGND _03874_ _03891_ keymem.prev_key0_reg\[104\] _03892_ sky130_fd_sc_hd__mux2_2
X_13064_ VGND VPWR _08577_ _07534_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_265_758 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_1044 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12015_ VGND VPWR VGND VPWR _07610_ keymem.key_mem\[7\]\[1\] _07611_ _07615_ _07617_
+ _07616_ sky130_fd_sc_hd__a2111o_2
X_17872_ VGND VPWR VPWR VGND _03836_ _03844_ keymem.prev_key0_reg\[82\] _03845_ sky130_fd_sc_hd__mux2_2
XFILLER_0_178_1157 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19611_ VGND VPWR _00598_ _05208_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_219_Right_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16823_ VGND VPWR _00053_ _02965_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_195_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_206_858 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19542_ VGND VPWR VPWR VGND _05151_ _04977_ keymem.key_mem\[12\]\[66\] _05172_ sky130_fd_sc_hd__mux2_2
X_13966_ VPWR VGND VGND VPWR _09432_ _09435_ _09436_ _09437_ _09438_ sky130_fd_sc_hd__and4b_2
X_16754_ VPWR VGND VPWR VGND _02902_ _02497_ _02898_ key[163] _02723_ _02903_ sky130_fd_sc_hd__a221o_2
XFILLER_0_205_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1346 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_92_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_152_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12917_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[75\] _07667_ keymem.key_mem\[7\]\[75\]
+ _07702_ _08445_ sky130_fd_sc_hd__a22o_2
XFILLER_0_156_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15705_ VPWR VGND _11161_ _11160_ keymem.prev_key0_reg\[16\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_19473_ VGND VPWR _05135_ _05092_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16685_ VGND VPWR _02839_ _02838_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13897_ VGND VPWR VGND VPWR _09369_ _09364_ _09363_ _09368_ _09367_ _09360_ sky130_fd_sc_hd__a32o_2
XFILLER_0_92_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_53_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18424_ VPWR VGND VPWR VGND _04312_ enc_block.round_key\[64\] _04311_ sky130_fd_sc_hd__or2_2
XFILLER_0_5_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15636_ VPWR VGND VPWR VGND _11094_ _11056_ sky130_fd_sc_hd__inv_2
X_12848_ VPWR VGND VPWR VGND _08382_ keymem.key_mem\[12\]\[68\] _07579_ keymem.key_mem\[4\]\[68\]
+ _07552_ _08383_ sky130_fd_sc_hd__a221o_2
XFILLER_0_29_624 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_56_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_61_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18355_ VPWR VGND VPWR VGND _04251_ _03996_ _04250_ sky130_fd_sc_hd__or2_2
X_15567_ VPWR VGND VPWR VGND _11026_ keymem.prev_key0_reg\[13\] sky130_fd_sc_hd__inv_2
X_12779_ VPWR VGND VPWR VGND _08320_ keymem.key_mem\[6\]\[61\] _07771_ keymem.key_mem\[10\]\[61\]
+ _07561_ _08321_ sky130_fd_sc_hd__a221o_2
X_14518_ VGND VPWR _09987_ _08935_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_124_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17306_ VGND VPWR VPWR VGND _03384_ keymem.key_mem\[14\]\[88\] _03401_ _03402_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_228_Right_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15498_ VGND VPWR VGND VPWR _10608_ _10575_ _10627_ _10498_ _10958_ sky130_fd_sc_hd__o22a_2
XFILLER_0_16_329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_638 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_18286_ VGND VPWR _04189_ _03950_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_43_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14449_ VGND VPWR VGND VPWR _09423_ _09330_ _09441_ _09355_ _09368_ _09918_ sky130_fd_sc_hd__o32a_2
X_17237_ VGND VPWR VPWR VGND _03296_ keymem.key_mem\[14\]\[81\] _03339_ _03340_ sky130_fd_sc_hd__mux2_2
XFILLER_0_265_1163 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_141_301 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_863 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_163_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_101_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17168_ VPWR VGND _03276_ _03278_ _03277_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_163_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_267 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_141_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16119_ VGND VPWR VGND VPWR _11236_ _11464_ _11380_ _11308_ _11573_ sky130_fd_sc_hd__o22a_2
XFILLER_0_229_906 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_60_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17099_ VPWR VGND VPWR VGND _03215_ _02497_ _09928_ key[195] _03211_ _03216_ sky130_fd_sc_hd__a221o_2
XFILLER_0_122_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_143_1_Right_744 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19809_ VGND VPWR _05314_ _05246_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_209_696 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_193_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22820_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[119\] _06860_ _06859_ _05073_ _02155_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_174_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_237_1276 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_56_1062 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22751_ VGND VPWR _02105_ _06841_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_71_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_21702_ VGND VPWR _01577_ _06320_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_17_1057 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_250_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25470_ VGND VPWR VPWR VGND clk _01963_ reset_n keymem.key_mem\[1\]\[55\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_66_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22682_ VGND VPWR VPWR VGND _06809_ keymem.key_mem\[0\]\[29\] _02812_ _06813_ sky130_fd_sc_hd__mux2_2
XFILLER_0_176_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_47_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24421_ VGND VPWR VPWR VGND clk _00914_ reset_n keymem.key_mem\[9\]\[30\] sky130_fd_sc_hd__dfrtp_2
X_21633_ VGND VPWR VPWR VGND _06275_ _02549_ keymem.key_mem\[4\]\[21\] _06284_ sky130_fd_sc_hd__mux2_2
XFILLER_0_191_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_605 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_142_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_627 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_69_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24352_ VGND VPWR VPWR VGND clk _00845_ reset_n keymem.key_mem\[10\]\[89\] sky130_fd_sc_hd__dfrtp_2
X_21564_ VGND VPWR _01513_ _06246_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_111_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_74_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23303_ VPWR VGND _07184_ enc_block.block_w1_reg\[9\] enc_block.block_w3_reg\[26\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_20515_ VGND VPWR VPWR VGND _05680_ _10835_ keymem.key_mem\[8\]\[10\] _05689_ sky130_fd_sc_hd__mux2_2
X_24283_ VGND VPWR VPWR VGND clk _00776_ reset_n keymem.key_mem\[10\]\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_7_595 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21495_ VGND VPWR _01480_ _06210_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_181_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23234_ VPWR VGND VPWR VGND _07122_ _07117_ _07120_ sky130_fd_sc_hd__or2_2
XFILLER_0_132_345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20446_ VGND VPWR VPWR VGND _05649_ _03533_ keymem.key_mem\[9\]\[106\] _05652_ sky130_fd_sc_hd__mux2_2
XFILLER_0_181_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_261_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23165_ VGND VPWR VGND VPWR _02293_ _07067_ _06888_ keymem.prev_key1_reg\[116\] sky130_fd_sc_hd__o21a_2
X_20377_ VGND VPWR VPWR VGND _05614_ _03268_ keymem.key_mem\[9\]\[73\] _05616_ sky130_fd_sc_hd__mux2_2
XFILLER_0_30_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_28_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22116_ VGND VPWR _01770_ _06541_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_219_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23096_ VGND VPWR VGND VPWR _03422_ _06928_ _03425_ _07024_ sky130_fd_sc_hd__a21o_2
XFILLER_0_100_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_237_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_961 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_100_286 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22047_ VGND VPWR _01737_ _06505_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_255_1310 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_215_622 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_243_942 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13820_ VPWR VGND VPWR VGND _09280_ _09291_ _09285_ _09275_ _09292_ sky130_fd_sc_hd__or4_2
X_25806_ keymem.prev_key1_reg\[122\] clk _02299_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_23998_ VGND VPWR VPWR VGND clk _00491_ reset_n keymem.key_mem\[13\]\[119\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_202_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13751_ VGND VPWR VGND VPWR _09223_ _09040_ _09058_ _09051_ _09057_ sky130_fd_sc_hd__a211o_2
X_25737_ keymem.prev_key1_reg\[53\] clk _02230_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_15_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22949_ VGND VPWR VPWR VGND _06914_ _06936_ keymem.prev_key1_reg\[31\] _06937_ sky130_fd_sc_hd__mux2_2
XFILLER_0_253_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12702_ VPWR VGND VPWR VGND _08250_ keymem.key_mem\[13\]\[54\] _07835_ keymem.key_mem\[4\]\[54\]
+ _07841_ _08251_ sky130_fd_sc_hd__a221o_2
X_16470_ VPWR VGND VPWR VGND _11514_ _11499_ _11529_ _11487_ _02631_ sky130_fd_sc_hd__or4_2
XFILLER_0_74_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13682_ VGND VPWR _09154_ _09072_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25668_ VGND VPWR VPWR VGND clk _02161_ reset_n keymem.key_mem\[0\]\[125\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15421_ VGND VPWR VGND VPWR _10528_ _10498_ _10882_ _10609_ sky130_fd_sc_hd__a21oi_2
X_12633_ VPWR VGND VPWR VGND _08188_ keymem.key_mem\[14\]\[47\] _07706_ keymem.key_mem\[2\]\[47\]
+ _07733_ _08189_ sky130_fd_sc_hd__a221o_2
X_24619_ VGND VPWR VPWR VGND clk _01112_ reset_n keymem.key_mem\[8\]\[100\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25599_ VGND VPWR VPWR VGND clk _02092_ reset_n keymem.key_mem\[0\]\[56\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_31_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15352_ VPWR VGND VGND VPWR _10785_ _10793_ _10813_ _10814_ sky130_fd_sc_hd__nor3_2
X_18140_ VPWR VGND _04055_ enc_block.block_w0_reg\[31\] enc_block.block_w0_reg\[30\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_12564_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[41\] _08125_ keymem.key_mem\[4\]\[41\]
+ _07693_ _08126_ sky130_fd_sc_hd__a22o_2
XFILLER_0_0_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14303_ VGND VPWR VGND VPWR _09386_ _09431_ _09564_ _09401_ _09773_ sky130_fd_sc_hd__o22a_2
X_18071_ VGND VPWR _03992_ _03949_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_108_386 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15283_ VGND VPWR VGND VPWR _08930_ key[137] _10745_ _10746_ sky130_fd_sc_hd__a21o_2
X_12495_ VGND VPWR VGND VPWR _08064_ _08008_ keymem.key_mem\[2\]\[34\] _08061_ _08063_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_227_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_800 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_660 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17022_ _02779_ _03146_ keymem.prev_key1_reg\[60\] _02780_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_14234_ VPWR VGND VGND VPWR _09140_ _09705_ _09082_ sky130_fd_sc_hd__nor2_2
XFILLER_0_145_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_33_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14165_ VGND VPWR VPWR VGND _09635_ _09549_ _09546_ _09636_ sky130_fd_sc_hd__mux2_2
XFILLER_0_145_1178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13116_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[95\] _07652_ keymem.key_mem\[8\]\[95\]
+ _08211_ _08624_ sky130_fd_sc_hd__a22o_2
XFILLER_0_237_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_260_1093 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14096_ VGND VPWR _09566_ _09397_ _09567_ _09564_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_18973_ VPWR VGND VPWR VGND _04806_ _04788_ _04805_ enc_block.block_w2_reg\[22\]
+ _04709_ _00362_ sky130_fd_sc_hd__a221o_2
XFILLER_0_81_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17924_ VGND VPWR _00239_ _03880_ VPWR VGND sky130_fd_sc_hd__buf_1
X_13047_ VGND VPWR VGND VPWR _07584_ keymem.key_mem\[14\]\[88\] _08559_ _08561_ _08562_
+ _08480_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_265_599 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_920 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17855_ VGND VPWR VGND VPWR _03304_ keymem.prev_key1_reg\[77\] _03833_ _03818_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_238_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_1_Left_382 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_245_290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_252_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_227_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16806_ VGND VPWR VGND VPWR _02949_ _02342_ _10384_ _10655_ _02950_ sky130_fd_sc_hd__a31o_2
X_17786_ VGND VPWR _00196_ _03785_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14998_ VGND VPWR _10462_ _10461_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_156_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19525_ VPWR VGND keymem.key_mem\[12\]\[58\] _05163_ _05158_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_88_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16737_ VGND VPWR VPWR VGND _10091_ key[162] keymem.prev_key1_reg\[34\] _02887_ sky130_fd_sc_hd__mux2_2
XFILLER_0_117_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13949_ VPWR VGND VPWR VGND _09261_ _09317_ _09314_ _09297_ _09421_ sky130_fd_sc_hd__or4_2
XFILLER_0_57_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_88_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_241_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_850 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_92_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19456_ VPWR VGND keymem.key_mem\[12\]\[26\] _05126_ _05116_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_53_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16668_ VPWR VGND VGND VPWR _02821_ _02820_ _10360_ _02818_ _02819_ _02822_ sky130_fd_sc_hd__a311o_2
XFILLER_0_134_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_158_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18407_ _04296_ _04298_ _04294_ _04297_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_118_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15619_ VPWR VGND VPWR VGND _11076_ _11077_ _10936_ _10991_ sky130_fd_sc_hd__or3b_2
XFILLER_0_201_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19387_ VGND VPWR VPWR VGND _05067_ _05085_ keymem.key_mem\[13\]\[125\] _05086_ sky130_fd_sc_hd__mux2_2
XFILLER_0_45_914 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16599_ VGND VPWR VGND VPWR _02747_ keymem.prev_key1_reg\[123\] _02756_ _02746_ sky130_fd_sc_hd__nand3_2
XFILLER_0_5_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18338_ VPWR VGND VPWR VGND _04236_ _03961_ _04234_ sky130_fd_sc_hd__or2_2
XFILLER_0_56_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18269_ VGND VPWR _04173_ enc_block.block_w1_reg\[17\] _04172_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_619 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_53_980 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20300_ VGND VPWR _00920_ _05575_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_163_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21280_ VGND VPWR VPWR VGND _06087_ _03567_ keymem.key_mem\[6\]\[112\] _06096_ sky130_fd_sc_hd__mux2_2
XFILLER_0_124_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_163_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20231_ VGND VPWR _00887_ _05539_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_188_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_64_1397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20162_ VGND VPWR VPWR VGND _05493_ _03499_ keymem.key_mem\[10\]\[101\] _05501_ sky130_fd_sc_hd__mux2_2
XFILLER_0_256_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24970_ VGND VPWR VPWR VGND clk _01463_ reset_n keymem.key_mem\[5\]\[67\] sky130_fd_sc_hd__dfrtp_2
X_20093_ VPWR VGND VGND VPWR _05465_ keymem.key_mem\[10\]\[68\] _05402_ sky130_fd_sc_hd__nand2_2
X_23921_ VGND VPWR VPWR VGND clk _00414_ reset_n keymem.key_mem\[13\]\[42\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_100_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_430 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_144_1_Right_745 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Right_2 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23852_ VGND VPWR VPWR VGND clk _00345_ reset_n enc_block.block_w2_reg\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_174_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22803_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[104\] _06858_ _06857_ _05041_ _02140_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_211_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23783_ VGND VPWR VPWR VGND clk _00276_ reset_n enc_block.block_w0_reg\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_75_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_135_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1227 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20995_ VGND VPWR _05945_ _05819_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_196_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_36_1444 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25522_ VGND VPWR VPWR VGND clk _02015_ reset_n keymem.key_mem\[1\]\[107\] sky130_fd_sc_hd__dfrtp_2
X_22734_ VGND VPWR VPWR VGND _06822_ keymem.key_mem\[0\]\[62\] _03173_ _06832_ sky130_fd_sc_hd__mux2_2
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25453_ VGND VPWR VPWR VGND clk _01946_ reset_n keymem.key_mem\[1\]\[38\] sky130_fd_sc_hd__dfrtp_2
X_22665_ VGND VPWR VPWR VGND _06798_ keymem.key_mem\[0\]\[21\] _02550_ _06804_ sky130_fd_sc_hd__mux2_2
XFILLER_0_149_297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24404_ VGND VPWR VPWR VGND clk _00897_ reset_n keymem.key_mem\[9\]\[13\] sky130_fd_sc_hd__dfrtp_2
X_21616_ VGND VPWR _06275_ _06262_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25384_ VGND VPWR VPWR VGND clk _01877_ reset_n keymem.key_mem\[2\]\[97\] sky130_fd_sc_hd__dfrtp_2
X_22596_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[108\] _06775_ _06774_ _05050_ _02016_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_168_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24335_ VGND VPWR VPWR VGND clk _00828_ reset_n keymem.key_mem\[10\]\[72\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_30_1087 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_21547_ VGND VPWR _01505_ _06237_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_181_1301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_248_1191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_146_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12280_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[16\] _07595_ keymem.key_mem\[6\]\[16\]
+ _07564_ _07867_ sky130_fd_sc_hd__a22o_2
X_24266_ VGND VPWR VPWR VGND clk _00759_ reset_n keymem.key_mem\[10\]\[3\] sky130_fd_sc_hd__dfrtp_2
X_21478_ VGND VPWR _01472_ _06201_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_82_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23217_ VGND VPWR _07106_ _03994_ _02306_ _07096_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_146_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20429_ VGND VPWR VPWR VGND _05638_ _03480_ keymem.key_mem\[9\]\[98\] _05643_ sky130_fd_sc_hd__mux2_2
X_24197_ VGND VPWR VPWR VGND clk _00690_ reset_n keymem.key_mem\[11\]\[62\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_181_1389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_685 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_219_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23148_ VGND VPWR VPWR VGND _07054_ _07057_ keymem.prev_key1_reg\[109\] _07058_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_180_1_Left_447 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_105_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15970_ VGND VPWR VGND VPWR _11426_ _11208_ _11228_ _11192_ _11288_ sky130_fd_sc_hd__and4_2
X_23079_ VGND VPWR VPWR VGND _06992_ _03354_ keymem.prev_key1_reg\[83\] _07015_ sky130_fd_sc_hd__mux2_2
XFILLER_0_41_1172 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_257_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14921_ VGND VPWR _10385_ keymem.prev_key0_reg\[8\] _10384_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_17640_ VGND VPWR VPWR VGND _03679_ key[134] keymem.prev_key1_reg\[6\] _03689_ sky130_fd_sc_hd__mux2_2
XFILLER_0_192_1430 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_463 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14852_ VGND VPWR _10317_ keymem.prev_key1_reg\[103\] _10316_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_153_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_794 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_192_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13803_ VGND VPWR VGND VPWR keymem.prev_key1_reg\[31\] _08969_ _09275_ _08964_ _09272_
+ _09274_ sky130_fd_sc_hd__a32oi_2
X_14783_ VGND VPWR VGND VPWR _09383_ _09352_ _10249_ _09323_ sky130_fd_sc_hd__a21oi_2
X_17571_ VGND VPWR VGND VPWR _03633_ _10838_ key[250] _03630_ _03632_ sky130_fd_sc_hd__a211o_2
XFILLER_0_93_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11995_ VPWR VGND VGND VPWR _07537_ _07598_ _07532_ sky130_fd_sc_hd__nor2_2
XFILLER_0_153_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19310_ VGND VPWR VPWR VGND _05025_ _05033_ keymem.key_mem\[13\]\[100\] _05034_ sky130_fd_sc_hd__mux2_2
X_13734_ VGND VPWR VGND VPWR _09206_ _09201_ _09199_ _09202_ _09205_ sky130_fd_sc_hd__a211o_2
X_16522_ VGND VPWR VGND VPWR _02679_ _02680_ _02682_ _02678_ sky130_fd_sc_hd__nand3_2
XFILLER_0_42_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_133_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19241_ VGND VPWR _00446_ _04990_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_196_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_16453_ VGND VPWR VGND VPWR _11295_ _11332_ _02614_ _11344_ sky130_fd_sc_hd__a21oi_2
X_13665_ VPWR VGND VPWR VGND _08963_ _09065_ _09051_ _09009_ _09137_ sky130_fd_sc_hd__or4_2
XFILLER_0_85_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_808 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15404_ VPWR VGND VPWR VGND _10864_ _10865_ _10862_ _10863_ sky130_fd_sc_hd__or3b_2
X_12616_ VGND VPWR enc_block.round_key\[45\] _08173_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16384_ VPWR VGND VPWR VGND _02547_ key[21] _11543_ sky130_fd_sc_hd__or2_2
X_19172_ VPWR VGND keymem.key_mem\[13\]\[47\] _04949_ _04915_ VPWR VGND sky130_fd_sc_hd__and2_2
X_13596_ VPWR VGND VPWR VGND _08963_ _09065_ _08971_ _09008_ _09068_ sky130_fd_sc_hd__or4_2
XFILLER_0_264_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15335_ VGND VPWR VPWR VGND _10430_ _10445_ _10424_ _10797_ sky130_fd_sc_hd__or3_2
X_18123_ VGND VPWR _04040_ _03950_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12547_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[39\] _07724_ keymem.key_mem\[1\]\[39\]
+ _07855_ _08111_ sky130_fd_sc_hd__a22o_2
XFILLER_0_170_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18054_ VGND VPWR VGND VPWR _03969_ _03951_ _03975_ _00274_ sky130_fd_sc_hd__a21o_2
X_15266_ _10677_ _10729_ keymem.round_ctr_reg\[0\] _10728_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_164_1543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12478_ VPWR VGND VPWR VGND _08047_ keymem.key_mem\[14\]\[33\] _08003_ keymem.key_mem\[6\]\[33\]
+ _07739_ _08048_ sky130_fd_sc_hd__a221o_2
XFILLER_0_41_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14217_ VGND VPWR VGND VPWR _09168_ _09136_ _09687_ _09688_ sky130_fd_sc_hd__a21o_2
XFILLER_0_125_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17005_ VGND VPWR VPWR VGND _03084_ keymem.key_mem\[14\]\[58\] _03130_ _03131_ sky130_fd_sc_hd__mux2_2
XFILLER_0_160_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15197_ VGND VPWR VGND VPWR _10661_ _10383_ _10382_ keylen _10660_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_21_140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_61_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14148_ VGND VPWR VGND VPWR _09434_ _09310_ _09440_ _09380_ _09247_ _09619_ sky130_fd_sc_hd__o32a_2
XFILLER_0_240_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_579 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_191_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_240_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14079_ VPWR VGND VGND VPWR _09304_ _09550_ _09319_ sky130_fd_sc_hd__nor2_2
X_18956_ VGND VPWR _04791_ enc_block.block_w1_reg\[5\] _04790_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_253_514 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17907_ VGND VPWR VPWR VGND _03792_ key[221] _03869_ _03868_ _03675_ sky130_fd_sc_hd__o211a_2
XFILLER_0_174_13 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18887_ VPWR VGND VPWR VGND _04729_ enc_block.block_w1_reg\[5\] enc_block.block_w1_reg\[6\]
+ sky130_fd_sc_hd__or2_2
XFILLER_0_207_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17838_ VGND VPWR VPWR VGND _03814_ _03821_ keymem.prev_key0_reg\[71\] _03822_ sky130_fd_sc_hd__mux2_2
XFILLER_0_171_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_233_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17769_ VGND VPWR _00189_ _03775_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_49_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19508_ VGND VPWR VPWR VGND _05151_ _04955_ keymem.key_mem\[12\]\[50\] _05154_ sky130_fd_sc_hd__mux2_2
X_20780_ VPWR VGND keymem.key_mem\[7\]\[5\] _05831_ _05830_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_14_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_499 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_212_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19439_ VPWR VGND keymem.key_mem\[12\]\[18\] _05117_ _05116_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_14_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_146_223 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_57_582 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22450_ VGND VPWR VPWR VGND _06715_ keymem.key_mem\[1\]\[19\] _02410_ _06719_ sky130_fd_sc_hd__mux2_2
XFILLER_0_91_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21401_ VGND VPWR VPWR VGND _06151_ _02955_ keymem.key_mem\[5\]\[40\] _06161_ sky130_fd_sc_hd__mux2_2
XFILLER_0_96_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22381_ VGND VPWR VPWR VGND _06680_ _03585_ keymem.key_mem\[2\]\[115\] _06682_ sky130_fd_sc_hd__mux2_2
XFILLER_0_5_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24120_ VGND VPWR VPWR VGND clk _00613_ reset_n keymem.key_mem\[12\]\[113\] sky130_fd_sc_hd__dfrtp_2
X_21332_ VGND VPWR VPWR VGND _06117_ _10369_ keymem.key_mem\[5\]\[7\] _06125_ sky130_fd_sc_hd__mux2_2
XFILLER_0_114_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_652 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24051_ VGND VPWR VPWR VGND clk _00544_ reset_n keymem.key_mem\[12\]\[44\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_114_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21263_ VGND VPWR _06087_ _05970_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_128_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23002_ VGND VPWR VPWR VGND _06960_ _06968_ keymem.prev_key1_reg\[52\] _06969_ sky130_fd_sc_hd__mux2_2
XFILLER_0_40_482 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20214_ VGND VPWR VPWR VGND _05388_ _03661_ keymem.key_mem\[10\]\[126\] _05528_ sky130_fd_sc_hd__mux2_2
XFILLER_0_25_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21194_ VGND VPWR VPWR VGND _06040_ _03251_ keymem.key_mem\[6\]\[71\] _06051_ sky130_fd_sc_hd__mux2_2
XFILLER_0_21_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_717 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_198_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20145_ VGND VPWR VPWR VGND _05482_ _03444_ keymem.key_mem\[10\]\[93\] _05492_ sky130_fd_sc_hd__mux2_2
XFILLER_0_99_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24953_ VGND VPWR VPWR VGND clk _01446_ reset_n keymem.key_mem\[5\]\[50\] sky130_fd_sc_hd__dfrtp_2
X_20076_ VGND VPWR VPWR VGND _05446_ _03150_ keymem.key_mem\[10\]\[60\] _05456_ sky130_fd_sc_hd__mux2_2
X_23904_ VGND VPWR VPWR VGND clk _00397_ reset_n keymem.key_mem\[13\]\[25\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_217_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24884_ VGND VPWR VPWR VGND clk _01377_ reset_n keymem.key_mem\[6\]\[109\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_169_304 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_145_1_Right_746 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23835_ VGND VPWR VPWR VGND clk _00328_ reset_n enc_block.block_w1_reg\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_139_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_197_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_36_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11780_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[25\] dec_new_block\[57\]
+ _07454_ sky130_fd_sc_hd__mux2_2
X_23766_ keymem.prev_key0_reg\[122\] clk _00263_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_20978_ VGND VPWR _01237_ _05936_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_71_1154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_135_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22717_ VGND VPWR VPWR VGND _06822_ keymem.key_mem\[0\]\[53\] _03083_ _06824_ sky130_fd_sc_hd__mux2_2
X_25505_ VGND VPWR VPWR VGND clk _01998_ reset_n keymem.key_mem\[1\]\[90\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_379 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23697_ keymem.prev_key0_reg\[53\] clk _00194_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_94_154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_211_1043 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_250_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13450_ VPWR VGND VGND VPWR _07376_ _00001_ _08923_ sky130_fd_sc_hd__nor2_2
X_25436_ VGND VPWR VPWR VGND clk _01929_ reset_n keymem.key_mem\[1\]\[21\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22648_ VGND VPWR VPWR VGND _06785_ keymem.key_mem\[0\]\[13\] _11040_ _06795_ sky130_fd_sc_hd__mux2_2
XFILLER_0_35_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_211_1098 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12401_ VGND VPWR VGND VPWR _07734_ keymem.key_mem\[4\]\[26\] _07975_ _07977_ _07978_
+ _07662_ sky130_fd_sc_hd__a2111o_2
X_25367_ VGND VPWR VPWR VGND clk _01860_ reset_n keymem.key_mem\[2\]\[80\] sky130_fd_sc_hd__dfrtp_2
X_13381_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[121\] _07861_ keymem.key_mem\[12\]\[121\]
+ _07787_ _08863_ sky130_fd_sc_hd__a22o_2
XFILLER_0_192_395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22579_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[94\] _06767_ _06766_ _05021_ _02002_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_90_360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1_1272 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15120_ VGND VPWR VPWR VGND _10463_ _10477_ _10500_ _10584_ sky130_fd_sc_hd__or3_2
XFILLER_0_51_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24318_ VGND VPWR VPWR VGND clk _00811_ reset_n keymem.key_mem\[10\]\[55\] sky130_fd_sc_hd__dfrtp_2
X_12332_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[20\] _07844_ keymem.key_mem\[4\]\[20\]
+ _07914_ _07915_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_438 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_105_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25298_ VGND VPWR VPWR VGND clk _01791_ reset_n keymem.key_mem\[2\]\[11\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_146_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15051_ VPWR VGND VGND VPWR _10500_ _10515_ _10514_ sky130_fd_sc_hd__nor2_2
XFILLER_0_267_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12263_ VPWR VGND VPWR VGND _07850_ keymem.key_mem\[6\]\[15\] _07657_ keymem.key_mem\[8\]\[15\]
+ _07655_ _07851_ sky130_fd_sc_hd__a221o_2
X_24249_ VGND VPWR VPWR VGND clk _00742_ reset_n keymem.key_mem\[11\]\[114\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_107_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14002_ VGND VPWR VPWR VGND _09331_ _09300_ _09319_ _09474_ sky130_fd_sc_hd__or3_2
XFILLER_0_47_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12194_ VGND VPWR _07787_ _07577_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_248_864 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18810_ VPWR VGND VGND VPWR _04660_ _04656_ _04658_ sky130_fd_sc_hd__nand2_2
XFILLER_0_43_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19790_ VGND VPWR _00681_ _05304_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_37_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18741_ VPWR VGND VPWR VGND _04596_ block[32] _04351_ enc_block.block_w1_reg\[0\]
+ _03954_ _04597_ sky130_fd_sc_hd__a221o_2
XFILLER_0_263_856 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15953_ _11266_ _11409_ _11263_ _11180_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_14904_ VGND VPWR VGND VPWR _10369_ _10324_ _10321_ _10326_ _10368_ sky130_fd_sc_hd__a211o_2
X_18672_ VPWR VGND VPWR VGND _04535_ _04459_ _04534_ enc_block.block_w1_reg\[24\]
+ _04424_ _00332_ sky130_fd_sc_hd__a221o_2
X_15884_ VPWR VGND VGND VPWR _11266_ _11340_ _11263_ sky130_fd_sc_hd__nor2_2
XFILLER_0_37_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17623_ VGND VPWR VGND VPWR _03670_ keymem.prev_key1_reg\[1\] _09547_ _03677_ sky130_fd_sc_hd__a21o_2
XFILLER_0_118_1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_153_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14835_ VPWR VGND VGND VPWR _09403_ _10300_ _09559_ sky130_fd_sc_hd__nor2_2
XFILLER_0_157_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17554_ VPWR VGND VGND VPWR _10287_ _03618_ key[248] sky130_fd_sc_hd__nor2_2
X_14766_ VPWR VGND VPWR VGND _09361_ _10231_ _09248_ _10063_ _10232_ sky130_fd_sc_hd__a22o_2
XFILLER_0_53_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11978_ VPWR VGND VGND VPWR _07543_ _07581_ _07531_ sky130_fd_sc_hd__nor2_2
XFILLER_0_114_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16505_ VPWR VGND VPWR VGND _11438_ _02665_ keymem.rcon_reg\[0\] _02498_ sky130_fd_sc_hd__or3b_2
X_13717_ VPWR VGND VGND VPWR _09189_ _09041_ _09086_ sky130_fd_sc_hd__nand2_2
X_14697_ VGND VPWR VGND VPWR _09177_ _09128_ _09146_ _09103_ _10164_ sky130_fd_sc_hd__o22a_2
X_17485_ VGND VPWR VPWR VGND _09730_ _11105_ key[239] _03558_ sky130_fd_sc_hd__mux2_2
XFILLER_0_6_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_316 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_85_187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19224_ VGND VPWR VGND VPWR _04980_ keymem.key_mem_we _03217_ _04968_ _00439_ sky130_fd_sc_hd__a31o_2
X_16436_ VGND VPWR VPWR VGND _11072_ _11089_ keymem.prev_key1_reg\[118\] _02598_ sky130_fd_sc_hd__or3_2
X_13648_ VPWR VGND VPWR VGND _08982_ _08997_ _08990_ _09001_ _09120_ sky130_fd_sc_hd__or4_2
XFILLER_0_128_267 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_89_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19155_ VGND VPWR VPWR VGND _04928_ _04937_ keymem.key_mem\[13\]\[41\] _04938_ sky130_fd_sc_hd__mux2_2
X_16367_ VGND VPWR VGND VPWR _11330_ _11352_ _02530_ _11311_ sky130_fd_sc_hd__a21oi_2
X_13579_ VGND VPWR _09051_ _09017_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18106_ VPWR VGND _04024_ enc_block.block_w0_reg\[28\] enc_block.block_w1_reg\[20\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_204_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_287 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15318_ VPWR VGND VPWR VGND _10778_ _10779_ _10780_ _10710_ _10777_ sky130_fd_sc_hd__or4b_2
X_16298_ VPWR VGND _02462_ keymem.prev_key0_reg\[84\] keymem.prev_key0_reg\[52\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
X_19086_ VGND VPWR VGND VPWR _04897_ keymem.key_mem_we _10977_ _04896_ _00384_ sky130_fd_sc_hd__a31o_2
XFILLER_0_78_11 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_164_1351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18037_ VGND VPWR _03959_ _03958_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15249_ VPWR VGND VPWR VGND _10710_ _10711_ _10712_ _10708_ _10709_ sky130_fd_sc_hd__or4b_2
XFILLER_0_151_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_26_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_164_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_188_2_Right_260 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_239_886 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_199_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19988_ VGND VPWR VPWR VGND _05400_ _02340_ keymem.key_mem\[10\]\[18\] _05410_ sky130_fd_sc_hd__mux2_2
XFILLER_0_226_536 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_185_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_96_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18939_ VPWR VGND VPWR VGND _04775_ block[51] _04744_ enc_block.block_w3_reg\[19\]
+ _04666_ _04776_ sky130_fd_sc_hd__a221o_2
XFILLER_0_253_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21950_ VGND VPWR VPWR VGND _06449_ _04935_ keymem.key_mem\[3\]\[40\] _06454_ sky130_fd_sc_hd__mux2_2
XFILLER_0_207_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20901_ VPWR VGND keymem.key_mem\[7\]\[61\] _05896_ _05886_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_178_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_178_112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_136_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21881_ VGND VPWR VGND VPWR _06416_ keymem.key_mem_we _10662_ _06404_ _01660_ sky130_fd_sc_hd__a31o_2
XFILLER_0_175_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_302 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23620_ VGND VPWR VPWR VGND clk _00121_ reset_n keymem.key_mem\[14\]\[109\] sky130_fd_sc_hd__dfrtp_2
X_20832_ VPWR VGND keymem.key_mem\[7\]\[29\] _05859_ _05856_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_136_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_72_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23551_ VGND VPWR VPWR VGND clk _00052_ reset_n keymem.key_mem\[14\]\[40\] sky130_fd_sc_hd__dfrtp_2
X_20763_ VPWR VGND VGND VPWR _05818_ _05819_ keymem.round_ctr_reg\[3\] sky130_fd_sc_hd__nor2_2
XFILLER_0_33_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22502_ VGND VPWR _06739_ _06695_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_91_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_23482_ VPWR VGND _07344_ enc_block.block_w1_reg\[13\] enc_block.block_w3_reg\[28\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_20694_ VGND VPWR _01107_ _05782_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_9_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25221_ VGND VPWR VPWR VGND clk _01714_ reset_n keymem.key_mem\[3\]\[62\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_247_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22433_ VGND VPWR _01918_ _06710_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_220_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_736 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25152_ VGND VPWR VPWR VGND clk _01645_ reset_n keymem.key_mem\[4\]\[121\] sky130_fd_sc_hd__dfrtp_2
X_22364_ VGND VPWR VPWR VGND _06669_ _03538_ keymem.key_mem\[2\]\[107\] _06673_ sky130_fd_sc_hd__mux2_2
XFILLER_0_66_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_606 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_24103_ VGND VPWR VPWR VGND clk _00596_ reset_n keymem.key_mem\[12\]\[96\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_182_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21315_ VPWR VGND VPWR VGND _06115_ _06114_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_112 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25083_ VGND VPWR VPWR VGND clk _01576_ reset_n keymem.key_mem\[4\]\[52\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_279 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_22295_ VPWR VGND VGND VPWR _06637_ keymem.key_mem\[2\]\[74\] _06567_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_196_Right_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_143_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_471 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24034_ VGND VPWR VPWR VGND clk _00527_ reset_n keymem.key_mem\[12\]\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_104_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21246_ VGND VPWR _01363_ _06078_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_229_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_143_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21177_ VGND VPWR _01330_ _06042_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_258_1533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20128_ VGND VPWR _00840_ _05483_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_245_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12950_ VGND VPWR VGND VPWR _08050_ keymem.key_mem\[7\]\[78\] _08471_ _08472_ _08475_
+ _08474_ sky130_fd_sc_hd__a2111o_2
X_20059_ VGND VPWR _00807_ _05447_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24936_ VGND VPWR VPWR VGND clk _01429_ reset_n keymem.key_mem\[5\]\[33\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_260_848 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11901_ VGND VPWR result[117] _07514_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12881_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[71\] _08124_ _08412_ _08408_ enc_block.round_key\[71\]
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_154_1531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24867_ VGND VPWR VPWR VGND clk _01360_ reset_n keymem.key_mem\[6\]\[92\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_146_1_Right_747 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_115_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11832_ VGND VPWR VPWR VGND encdec enc_block.block_w1_reg\[19\] dec_new_block\[83\]
+ _07480_ sky130_fd_sc_hd__mux2_2
XFILLER_0_240_572 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14620_ VGND VPWR _10088_ keymem.prev_key1_reg\[100\] _10087_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_154_1575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23818_ VGND VPWR VPWR VGND clk _00311_ reset_n enc_block.block_w1_reg\[3\] sky130_fd_sc_hd__dfrtp_2
X_24798_ VGND VPWR VPWR VGND clk _01291_ reset_n keymem.key_mem\[6\]\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_90_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14551_ VPWR VGND VPWR VGND _10019_ _09185_ sky130_fd_sc_hd__inv_2
X_11763_ VGND VPWR result[48] _07445_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_230_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23749_ keymem.prev_key0_reg\[105\] clk _00246_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_3_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13502_ enc_block.sword_ctr_reg\[1\] _08974_ enc_block.sword_ctr_reg\[0\] enc_block.block_w3_reg\[7\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_51_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14482_ VPWR VGND VPWR VGND _09950_ _09951_ _09180_ _09813_ sky130_fd_sc_hd__or3b_2
X_17270_ VGND VPWR VGND VPWR _03368_ _03367_ _10386_ _03369_ sky130_fd_sc_hd__a21o_2
XFILLER_0_230_1485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11694_ VGND VPWR VPWR VGND encdec enc_block.block_w3_reg\[14\] dec_new_block\[14\]
+ _07411_ sky130_fd_sc_hd__mux2_2
X_16221_ VPWR VGND VGND VPWR _11527_ _02386_ _11314_ sky130_fd_sc_hd__nor2_2
X_13433_ VGND VPWR VGND VPWR _08910_ _08096_ keymem.key_mem\[5\]\[126\] _08907_ _08909_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_187_1362 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_265_1537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25419_ VGND VPWR VPWR VGND clk _01912_ reset_n keymem.key_mem\[1\]\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_130_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16152_ VGND VPWR VGND VPWR _11372_ _11332_ _11239_ _11606_ sky130_fd_sc_hd__a21o_2
X_13364_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[119\] _08027_ _08847_ _08843_ _08848_
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_180_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_63_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_124_1_Left_391 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15103_ VPWR VGND VGND VPWR _10566_ _10567_ _10565_ sky130_fd_sc_hd__nor2_2
X_12315_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[19\] _07702_ keymem.key_mem\[9\]\[19\]
+ _07716_ _07899_ sky130_fd_sc_hd__a22o_2
X_16083_ VGND VPWR VGND VPWR _11537_ _11535_ _11538_ _11536_ sky130_fd_sc_hd__nand3_2
XFILLER_0_133_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13295_ VGND VPWR enc_block.round_key\[112\] _08785_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_161_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15034_ VGND VPWR _10498_ _10497_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19911_ VGND VPWR _00739_ _05367_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12246_ VGND VPWR _07835_ _07834_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_122_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19842_ VGND VPWR _00706_ _05331_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12177_ VGND VPWR _07771_ _07564_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_236_834 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_202_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_536 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_200_Right_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_257_1021 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19773_ VGND VPWR _00673_ _05295_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16985_ VPWR VGND VPWR VGND _03112_ key[57] _09719_ sky130_fd_sc_hd__or2_2
XFILLER_0_262_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18724_ VPWR VGND _04582_ _04581_ enc_block.round_key\[94\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15936_ VPWR VGND VGND VPWR _11278_ _11392_ _11391_ sky130_fd_sc_hd__nor2_2
XFILLER_0_64_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18655_ VPWR VGND VGND VPWR _04512_ _04521_ _04223_ sky130_fd_sc_hd__nor2_2
X_15867_ VGND VPWR _11323_ _11222_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_59_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17606_ VPWR VGND VGND VPWR _03663_ _03240_ _02847_ sky130_fd_sc_hd__nand2_2
XFILLER_0_154_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14818_ VGND VPWR _10284_ _10283_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18586_ VGND VPWR _04459_ _03950_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15798_ VGND VPWR VGND VPWR _11253_ _11246_ _11250_ _11219_ _11254_ sky130_fd_sc_hd__a31o_2
XFILLER_0_118_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17537_ VPWR VGND VPWR VGND _03603_ key[118] _11543_ sky130_fd_sc_hd__or2_2
XFILLER_0_15_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14749_ VPWR VGND VGND VPWR _10199_ _10204_ _10209_ _10214_ _10215_ sky130_fd_sc_hd__and4b_2
XFILLER_0_58_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_699 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_171_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17468_ VGND VPWR VPWR VGND _03534_ keymem.key_mem\[14\]\[108\] _03543_ _03544_ sky130_fd_sc_hd__mux2_2
XFILLER_0_229_1101 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_116_204 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19207_ VGND VPWR VGND VPWR _04970_ keymem.key_mem_we _03150_ _04968_ _00432_ sky130_fd_sc_hd__a31o_2
X_16419_ VGND VPWR VPWR VGND _11278_ _11308_ _11477_ _02581_ sky130_fd_sc_hd__or3_2
XFILLER_0_89_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17399_ VPWR VGND _02496_ _03484_ _03483_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_229_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_27_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_171_354 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19138_ VGND VPWR VGND VPWR _04926_ keymem.key_mem_we _02904_ _04924_ _00407_ sky130_fd_sc_hd__a31o_2
XFILLER_0_42_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19069_ VGND VPWR _04887_ _04879_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_2_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21100_ VGND VPWR VPWR VGND _05996_ _02742_ keymem.key_mem\[6\]\[26\] _06002_ sky130_fd_sc_hd__mux2_2
XFILLER_0_164_1192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_203_1318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22080_ VGND VPWR _01753_ _06522_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_11_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21031_ VGND VPWR VPWR VGND _05956_ _05081_ keymem.key_mem\[7\]\[123\] _05964_ sky130_fd_sc_hd__mux2_2
XFILLER_0_59_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1186 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_10_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_189_2_Right_261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_201_1053 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_96_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_242_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_199_719 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_25770_ keymem.prev_key1_reg\[86\] clk _02263_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_22982_ VGND VPWR VPWR VGND _06914_ _06956_ keymem.prev_key1_reg\[44\] _06957_ sky130_fd_sc_hd__mux2_2
XFILLER_0_254_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_198_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24721_ VGND VPWR VPWR VGND clk _01214_ reset_n keymem.key_mem\[7\]\[74\] sky130_fd_sc_hd__dfrtp_2
X_21933_ VGND VPWR _01684_ _06444_ VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_168_2_Left_639 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_210_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_250_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24652_ VGND VPWR VPWR VGND clk _01145_ reset_n keymem.key_mem\[7\]\[5\] sky130_fd_sc_hd__dfrtp_2
X_21864_ VGND VPWR VGND VPWR _06407_ keymem.key_mem_we _09537_ _06404_ _01652_ sky130_fd_sc_hd__a31o_2
XFILLER_0_136_1283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23603_ VGND VPWR VPWR VGND clk _00104_ reset_n keymem.key_mem\[14\]\[92\] sky130_fd_sc_hd__dfrtp_2
X_20815_ VGND VPWR VGND VPWR _05849_ keymem.key_mem_we _02550_ _05838_ _01161_ sky130_fd_sc_hd__a31o_2
X_24583_ VGND VPWR VPWR VGND clk _01076_ reset_n keymem.key_mem\[8\]\[64\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21795_ VGND VPWR VPWR VGND _06366_ _03480_ keymem.key_mem\[4\]\[98\] _06369_ sky130_fd_sc_hd__mux2_2
XFILLER_0_166_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_1_Right_671 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_64_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23534_ VGND VPWR VPWR VGND clk _00035_ reset_n keymem.key_mem\[14\]\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_64_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20746_ VGND VPWR VPWR VGND _05805_ _03620_ keymem.key_mem\[8\]\[120\] _05810_ sky130_fd_sc_hd__mux2_2
XFILLER_0_9_251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_231_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23465_ VPWR VGND VGND VPWR _07329_ _07117_ _07328_ sky130_fd_sc_hd__nand2_2
X_20677_ VGND VPWR VPWR VGND _05772_ _03392_ keymem.key_mem\[8\]\[87\] _05774_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25204_ VGND VPWR VPWR VGND clk _01697_ reset_n keymem.key_mem\[3\]\[45\] sky130_fd_sc_hd__dfrtp_2
X_22416_ VGND VPWR _01911_ _06700_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23396_ VPWR VGND VPWR VGND _07268_ _07265_ _07267_ sky130_fd_sc_hd__or2_2
X_25135_ VGND VPWR VPWR VGND clk _01628_ reset_n keymem.key_mem\[4\]\[104\] sky130_fd_sc_hd__dfrtp_2
X_22347_ VGND VPWR VPWR VGND _06658_ _03485_ keymem.key_mem\[2\]\[99\] _06664_ sky130_fd_sc_hd__mux2_2
X_12100_ VGND VPWR _07698_ _07697_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_108_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13080_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[91\] _08391_ keymem.key_mem\[14\]\[91\]
+ _07632_ _08592_ sky130_fd_sc_hd__a22o_2
X_25066_ VGND VPWR VPWR VGND clk _01559_ reset_n keymem.key_mem\[4\]\[35\] sky130_fd_sc_hd__dfrtp_2
X_22278_ VGND VPWR VPWR VGND _06622_ _03209_ keymem.key_mem\[2\]\[66\] _06628_ sky130_fd_sc_hd__mux2_2
XFILLER_0_104_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12031_ VGND VPWR _07632_ _07582_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24017_ VGND VPWR VPWR VGND clk _00510_ reset_n keymem.key_mem\[12\]\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_44_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21229_ VGND VPWR _01355_ _06069_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_16770_ VGND VPWR VPWR VGND _10144_ _02916_ keymem.prev_key1_reg\[37\] _02917_ sky130_fd_sc_hd__mux2_2
XFILLER_0_258_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13982_ VGND VPWR VGND VPWR _09454_ _09448_ _09447_ _09451_ _09453_ sky130_fd_sc_hd__a211o_2
XFILLER_0_254_1249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15721_ VGND VPWR VGND VPWR enc_block.block_w2_reg\[17\] _09269_ _10387_ _11175_
+ _11177_ _11176_ sky130_fd_sc_hd__a2111o_2
X_12933_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[77\] _07984_ keymem.key_mem\[1\]\[77\]
+ _07969_ _08459_ sky130_fd_sc_hd__a22o_2
X_24919_ VGND VPWR VPWR VGND clk _01412_ reset_n keymem.key_mem\[5\]\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_1144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_18440_ VPWR VGND _04327_ _04326_ enc_block.round_key\[65\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_217_1071 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_87_238 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15652_ VGND VPWR _11109_ _09987_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_115_1323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_892 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12864_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[70\] _07659_ keymem.key_mem\[10\]\[70\]
+ _08193_ _08397_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_147_1_Right_748 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14603_ VGND VPWR VGND VPWR _09564_ _09353_ _10071_ _09411_ sky130_fd_sc_hd__a21oi_2
X_18371_ VGND VPWR _04266_ _04148_ VPWR VGND sky130_fd_sc_hd__buf_1
X_11815_ VGND VPWR result[74] _07471_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_115_1367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12795_ VPWR VGND VPWR VGND _08334_ keymem.key_mem\[3\]\[63\] _07844_ keymem.key_mem\[9\]\[63\]
+ _07738_ _08335_ sky130_fd_sc_hd__a221o_2
XFILLER_0_200_244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15583_ VGND VPWR VPWR VGND _11041_ keymem.key_mem\[14\]\[13\] _11040_ _11042_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_636 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_261_Right_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17322_ VGND VPWR VPWR VGND _03414_ _02691_ _03416_ _09722_ _03415_ sky130_fd_sc_hd__o211a_2
XFILLER_0_12_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11746_ VGND VPWR VPWR VGND encdec enc_block.block_w2_reg\[8\] dec_new_block\[40\]
+ _07437_ sky130_fd_sc_hd__mux2_2
X_14534_ VPWR VGND VPWR VGND _09841_ _10001_ _09997_ _09234_ _10002_ sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_1_Left_269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_850 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17253_ VGND VPWR VGND VPWR _03354_ _03351_ _03350_ _09534_ _03353_ _03349_ sky130_fd_sc_hd__a32o_2
XFILLER_0_138_395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14465_ VPWR VGND _09934_ _09933_ keymem.prev_key0_reg\[3\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_11677_ VGND VPWR result[5] _07402_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_153_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_265_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_917 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16204_ VGND VPWR VGND VPWR _11380_ _11375_ _11386_ _11473_ _02369_ sky130_fd_sc_hd__o22a_2
XFILLER_0_187_1192 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13416_ VPWR VGND VPWR VGND keymem.key_mem\[14\]\[125\] _07782_ keymem.key_mem\[10\]\[125\]
+ _07785_ _08894_ sky130_fd_sc_hd__a22o_2
XFILLER_0_3_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14396_ VGND VPWR _00014_ _09865_ VPWR VGND sky130_fd_sc_hd__buf_1
X_17184_ VGND VPWR _02866_ key[76] _03292_ _03029_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_221_83 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_10_1085 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_555 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_184 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16135_ VGND VPWR VGND VPWR _11572_ _11589_ _11583_ _11588_ _11577_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_45_1104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13347_ VGND VPWR VGND VPWR _08832_ _07841_ keymem.key_mem\[4\]\[118\] _08831_ _08020_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_224_1031 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_59_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16066_ _11230_ _11521_ _11391_ _11291_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_13278_ VPWR VGND VPWR VGND keymem.key_mem\[3\]\[111\] _07843_ keymem.key_mem\[2\]\[111\]
+ _07697_ _08770_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15017_ VGND VPWR VPWR VGND _10453_ _10409_ _10439_ _10481_ sky130_fd_sc_hd__or3_2
XFILLER_0_249_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12229_ VPWR VGND VPWR VGND _07819_ keymem.key_mem\[6\]\[12\] _07818_ keymem.key_mem\[9\]\[12\]
+ _07705_ _07820_ sky130_fd_sc_hd__a221o_2
XFILLER_0_209_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_202_1340 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_97_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19825_ VGND VPWR _00698_ _05322_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_209_867 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_97_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19756_ VGND VPWR _00665_ _05286_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_237_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16968_ VGND VPWR VGND VPWR _03096_ _03097_ _02655_ _02654_ sky130_fd_sc_hd__o21bai_2
X_18707_ VPWR VGND _04567_ _04566_ enc_block.round_key\[92\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_237_1469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15919_ VGND VPWR _11375_ _11307_ VPWR VGND sky130_fd_sc_hd__buf_1
X_19687_ VGND VPWR _00632_ _05250_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16899_ VPWR VGND VPWR VGND _03034_ _03031_ _03028_ key[176] _03027_ _03035_ sky130_fd_sc_hd__a221o_2
XFILLER_0_155_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18638_ VGND VPWR _04505_ _04103_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_91_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18569_ VGND VPWR _04443_ enc_block.block_w2_reg\[22\] enc_block.block_w1_reg\[30\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_496 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20600_ VGND VPWR _01062_ _05733_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21580_ VGND VPWR _01521_ _06254_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_46_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_129_362 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_850 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20531_ VGND VPWR _01029_ _05697_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_7_755 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_209_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_144_343 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_248_1565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_691 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23250_ VPWR VGND _07137_ _07136_ enc_block.round_key\[4\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_6_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20462_ VGND VPWR _05660_ _05533_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_244_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_1_Right_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22201_ VGND VPWR _01809_ _06587_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_259_712 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23181_ VGND VPWR VGND VPWR _03636_ _03635_ _03639_ _07077_ sky130_fd_sc_hd__a21o_2
XFILLER_0_43_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20393_ VGND VPWR VPWR VGND _05614_ _03339_ keymem.key_mem\[9\]\[81\] _05624_ sky130_fd_sc_hd__mux2_2
XFILLER_0_30_536 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_105_1503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22132_ VGND VPWR _01778_ _06549_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_144_1563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22063_ VGND VPWR VGND VPWR _06513_ keymem.key_mem_we _03444_ _06498_ _01745_ sky130_fd_sc_hd__a31o_2
X_21014_ VGND VPWR VPWR VGND _05945_ _05064_ keymem.key_mem\[7\]\[115\] _05955_ sky130_fd_sc_hd__mux2_2
XFILLER_0_226_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25822_ VGND VPWR VPWR VGND clk _02315_ reset_n enc_block.block_w3_reg\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_254_472 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_255_1525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22965_ VGND VPWR VPWR VGND _06914_ _06946_ keymem.prev_key1_reg\[37\] _06947_ sky130_fd_sc_hd__mux2_2
X_25753_ keymem.prev_key1_reg\[69\] clk _02246_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_24704_ VGND VPWR VPWR VGND clk _01197_ reset_n keymem.key_mem\[7\]\[57\] sky130_fd_sc_hd__dfrtp_2
X_21916_ VGND VPWR VGND VPWR _06435_ keymem.key_mem_we _02689_ _06432_ _01676_ sky130_fd_sc_hd__a31o_2
XFILLER_0_69_249 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22896_ VGND VPWR VGND VPWR _02188_ _06903_ _06882_ keymem.prev_key1_reg\[11\] sky130_fd_sc_hd__o21a_2
X_25684_ keymem.prev_key1_reg\[0\] clk _02177_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_222_391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_112_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24635_ VGND VPWR VPWR VGND clk _01128_ reset_n keymem.key_mem\[8\]\[116\] sky130_fd_sc_hd__dfrtp_2
X_21847_ VGND VPWR VPWR VGND _06388_ _03640_ keymem.key_mem\[4\]\[123\] _06396_ sky130_fd_sc_hd__mux2_2
XFILLER_0_214_1288 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_139_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_37_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_249_1307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24566_ VGND VPWR VPWR VGND clk _01059_ reset_n keymem.key_mem\[8\]\[47\] sky130_fd_sc_hd__dfrtp_2
X_12580_ VPWR VGND VPWR VGND keymem.key_mem\[9\]\[42\] _07612_ keymem.key_mem\[4\]\[42\]
+ _07692_ _08141_ sky130_fd_sc_hd__a22o_2
XFILLER_0_194_265 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_38_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_1_Right_672 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_249_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21778_ VGND VPWR VPWR VGND _06355_ _03417_ keymem.key_mem\[4\]\[90\] _06360_ sky130_fd_sc_hd__mux2_2
X_23517_ VGND VPWR VPWR VGND clk _00018_ reset_n keymem.key_mem\[14\]\[6\] sky130_fd_sc_hd__dfrtp_2
X_20729_ VGND VPWR VPWR VGND _05794_ _03567_ keymem.key_mem\[8\]\[112\] _05801_ sky130_fd_sc_hd__mux2_2
X_24497_ VGND VPWR VPWR VGND clk _00990_ reset_n keymem.key_mem\[9\]\[106\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_110_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14250_ VGND VPWR _09721_ _09512_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23448_ VGND VPWR VPWR VGND _07312_ _07247_ _07314_ _03982_ _07313_ sky130_fd_sc_hd__o211a_2
XFILLER_0_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13201_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[103\] _08193_ keymem.key_mem\[12\]\[103\]
+ _07620_ _08701_ sky130_fd_sc_hd__a22o_2
X_14181_ VPWR VGND VGND VPWR _09646_ _09127_ _09652_ _09154_ _09102_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_184_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_909 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_23379_ VPWR VGND VPWR VGND _07252_ block[17] _04837_ enc_block.block_w0_reg\[17\]
+ _04504_ _07253_ sky130_fd_sc_hd__a221o_2
XFILLER_0_249_211 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_61_694 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13132_ VPWR VGND VPWR VGND _08638_ keymem.key_mem\[11\]\[96\] _07912_ keymem.key_mem\[1\]\[96\]
+ _07969_ _08639_ sky130_fd_sc_hd__a221o_2
X_25118_ VGND VPWR VPWR VGND clk _01611_ reset_n keymem.key_mem\[4\]\[87\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_81_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_108_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_237_417 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_29_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17940_ VGND VPWR VGND VPWR _03515_ keymem.prev_key1_reg\[104\] _03891_ _03818_ sky130_fd_sc_hd__a21bo_2
X_13063_ VGND VPWR enc_block.round_key\[89\] _08576_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_221_1248 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25049_ VGND VPWR VPWR VGND clk _01542_ reset_n keymem.key_mem\[4\]\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_267_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_428 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12014_ VGND VPWR _07616_ _07572_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_79_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17871_ VGND VPWR VPWR VGND _03812_ key[210] keymem.prev_key1_reg\[82\] _03844_ sky130_fd_sc_hd__mux2_2
XFILLER_0_40_1056 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19610_ VGND VPWR VPWR VGND _05205_ _05029_ keymem.key_mem\[12\]\[98\] _05208_ sky130_fd_sc_hd__mux2_2
XFILLER_0_79_1255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16822_ VGND VPWR VPWR VGND _02884_ keymem.key_mem\[14\]\[41\] _02964_ _02965_ sky130_fd_sc_hd__mux2_2
XFILLER_0_218_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19541_ VGND VPWR _00565_ _05171_ VPWR VGND sky130_fd_sc_hd__buf_1
X_16753_ VGND VPWR VGND VPWR _02899_ _09933_ _02902_ _02901_ sky130_fd_sc_hd__a21oi_2
X_13965_ VPWR VGND VGND VPWR _09437_ _09319_ _09331_ sky130_fd_sc_hd__nand2_2
XFILLER_0_221_818 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15704_ VPWR VGND _11160_ keymem.prev_key0_reg\[80\] keymem.prev_key0_reg\[48\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
X_19472_ VGND VPWR _00533_ _05134_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12916_ VPWR VGND VPWR VGND keymem.key_mem\[4\]\[75\] _07734_ keymem.key_mem\[2\]\[75\]
+ _08131_ _08444_ sky130_fd_sc_hd__a22o_2
XFILLER_0_220_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16684_ VPWR VGND VPWR VGND _02837_ _02677_ _02827_ key[158] _02723_ _02838_ sky130_fd_sc_hd__a221o_2
X_13896_ VGND VPWR _09368_ _09362_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18423_ VPWR VGND VPWR VGND _04310_ block[64] _03980_ enc_block.block_w0_reg\[0\]
+ _03978_ _04311_ sky130_fd_sc_hd__a221o_2
XFILLER_0_57_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15635_ VPWR VGND VGND VPWR _11092_ _11093_ _10386_ sky130_fd_sc_hd__nor2_2
XFILLER_0_185_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12847_ VPWR VGND VPWR VGND keymem.key_mem\[5\]\[68\] _07596_ keymem.key_mem\[7\]\[68\]
+ _07609_ _08382_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_148_1_Right_749 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_8_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18354_ VGND VPWR _04250_ enc_block.block_w3_reg\[2\] _03985_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15566_ VGND VPWR VGND VPWR _11022_ _11021_ _11023_ _11025_ sky130_fd_sc_hd__a21o_2
X_12778_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[61\] _07608_ keymem.key_mem\[9\]\[61\]
+ _07591_ _08320_ sky130_fd_sc_hd__a22o_2
XFILLER_0_267_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17305_ VPWR VGND VPWR VGND _03400_ _10902_ _03398_ key[216] _03366_ _03401_ sky130_fd_sc_hd__a221o_2
XFILLER_0_56_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14517_ VGND VPWR VPWR VGND _09934_ _09985_ _09932_ _09986_ sky130_fd_sc_hd__or3_2
X_18285_ VPWR VGND _04188_ _04187_ enc_block.round_key\[115\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_11729_ VGND VPWR result[31] _07428_ VPWR VGND sky130_fd_sc_hd__buf_1
X_15497_ VGND VPWR VGND VPWR _10547_ _10583_ _10515_ _10628_ _10646_ _10957_ sky130_fd_sc_hd__o32a_2
XFILLER_0_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_831 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17236_ VPWR VGND VPWR VGND _03338_ _03336_ _03335_ key[209] _03027_ _03339_ sky130_fd_sc_hd__a221o_2
XFILLER_0_117_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14448_ VPWR VGND VPWR VGND _09914_ _09916_ _09915_ _09913_ _09917_ sky130_fd_sc_hd__or4_2
XFILLER_0_43_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_725 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_875 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17167_ VPWR VGND VGND VPWR _03277_ key[202] _08930_ sky130_fd_sc_hd__nand2_2
XFILLER_0_25_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14379_ VPWR VGND VPWR VGND _09848_ _09849_ _09846_ _09847_ sky130_fd_sc_hd__or3b_2
X_16118_ VPWR VGND VPWR VGND _11570_ _11571_ _11572_ _11563_ _11568_ sky130_fd_sc_hd__or4b_2
X_17098_ VGND VPWR VPWR VGND _03212_ keymem.prev_key0_reg\[67\] _03215_ _03214_ _03213_
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_0_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16049_ VPWR VGND VGND VPWR _11314_ _11504_ _11205_ sky130_fd_sc_hd__nor2_2
XFILLER_0_256_737 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_122_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_19808_ VGND VPWR _00690_ _05313_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_19_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_792 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_263_291 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_193_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_100_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_223_144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19739_ VGND VPWR _00657_ _05277_ VPWR VGND sky130_fd_sc_hd__buf_1
X_22750_ VGND VPWR VPWR VGND _06833_ keymem.key_mem\[0\]\[69\] _03235_ _06841_ sky130_fd_sc_hd__mux2_2
XFILLER_0_35_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21701_ VGND VPWR VPWR VGND _06319_ _03082_ keymem.key_mem\[4\]\[53\] _06320_ sky130_fd_sc_hd__mux2_2
X_22681_ VGND VPWR _02064_ _06812_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_250_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24420_ VGND VPWR VPWR VGND clk _00913_ reset_n keymem.key_mem\[9\]\[29\] sky130_fd_sc_hd__dfrtp_2
X_21632_ VGND VPWR _01544_ _06283_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_47_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_142_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24351_ VGND VPWR VPWR VGND clk _00844_ reset_n keymem.key_mem\[10\]\[88\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_129_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21563_ VGND VPWR VPWR VGND _06242_ _03600_ keymem.key_mem\[5\]\[117\] _06246_ sky130_fd_sc_hd__mux2_2
XFILLER_0_63_937 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_69_1435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23302_ VGND VPWR _07183_ _04086_ _02314_ _07096_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_191_268 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_20514_ VGND VPWR _01021_ _05688_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_248_1373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24282_ VGND VPWR VPWR VGND clk _00775_ reset_n keymem.key_mem\[10\]\[19\] sky130_fd_sc_hd__dfrtp_2
X_21494_ VGND VPWR VPWR VGND _06209_ _03364_ keymem.key_mem\[5\]\[84\] _06210_ sky130_fd_sc_hd__mux2_2
XFILLER_0_27_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_69_1479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23233_ VPWR VGND VGND VPWR _07121_ _07117_ _07120_ sky130_fd_sc_hd__nand2_2
XFILLER_0_181_1527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20445_ VGND VPWR _00989_ _05651_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_132_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23164_ VGND VPWR VGND VPWR _07067_ _03588_ _06890_ _03591_ _07011_ sky130_fd_sc_hd__a211o_2
XFILLER_0_105_1311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20376_ VGND VPWR _00956_ _05615_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_109_1491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22115_ VGND VPWR VPWR VGND _06538_ _05071_ keymem.key_mem\[3\]\[118\] _06541_ sky130_fd_sc_hd__mux2_2
XFILLER_0_100_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23095_ VGND VPWR _02267_ _07023_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_179_1423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22046_ VGND VPWR VPWR VGND _06494_ _05008_ keymem.key_mem\[3\]\[85\] _06505_ sky130_fd_sc_hd__mux2_2
XFILLER_0_237_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_133 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25805_ keymem.prev_key1_reg\[121\] clk _02298_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_199_346 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23997_ VGND VPWR VPWR VGND clk _00490_ reset_n keymem.key_mem\[13\]\[118\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_253_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13750_ VGND VPWR _09222_ _09121_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25736_ keymem.prev_key1_reg\[52\] clk _02229_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_202_328 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22948_ VGND VPWR VGND VPWR _02851_ _06928_ _02860_ _06936_ sky130_fd_sc_hd__a21o_2
XPHY_EDGE_ROW_101_2_Left_572 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12701_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[54\] _07562_ keymem.key_mem\[1\]\[54\]
+ _07558_ _08250_ sky130_fd_sc_hd__a22o_2
XFILLER_0_211_851 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_1147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13681_ VGND VPWR _09153_ _09029_ VPWR VGND sky130_fd_sc_hd__buf_1
X_25667_ VGND VPWR VPWR VGND clk _02160_ reset_n keymem.key_mem\[0\]\[124\] sky130_fd_sc_hd__dfrtp_2
X_22879_ VGND VPWR VGND VPWR _02181_ _06893_ _06882_ keymem.prev_key1_reg\[4\] sky130_fd_sc_hd__o21a_2
XFILLER_0_13_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15420_ VPWR VGND VPWR VGND _10878_ _10517_ _10879_ _10880_ _10881_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_17_1581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12632_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[47\] _07674_ keymem.key_mem\[4\]\[47\]
+ _07692_ _08188_ sky130_fd_sc_hd__a22o_2
X_24618_ VGND VPWR VPWR VGND clk _01111_ reset_n keymem.key_mem\[8\]\[99\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_167_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_25598_ VGND VPWR VPWR VGND clk _02091_ reset_n keymem.key_mem\[0\]\[55\] sky130_fd_sc_hd__dfrtp_2
X_15351_ VPWR VGND VPWR VGND _10801_ _10812_ _10806_ _10795_ _10813_ sky130_fd_sc_hd__or4_2
XFILLER_0_108_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12563_ VGND VPWR _08125_ _07694_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_25_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_1_Right_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24549_ VGND VPWR VPWR VGND clk _01042_ reset_n keymem.key_mem\[8\]\[30\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_87_1535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14302_ VGND VPWR VPWR VGND _09367_ _09626_ _09295_ _09772_ sky130_fd_sc_hd__or3_2
X_18070_ VPWR VGND _03991_ _03990_ enc_block.round_key\[97\] VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_0_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_123_302 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12494_ VPWR VGND VPWR VGND _08062_ keymem.key_mem\[14\]\[34\] _07706_ keymem.key_mem\[11\]\[34\]
+ _07902_ _08063_ sky130_fd_sc_hd__a221o_2
X_15282_ VPWR VGND VGND VPWR _10734_ _10736_ _10745_ _10744_ _10743_ sky130_fd_sc_hd__o22ai_2
XPHY_EDGE_ROW_152_1_Left_419 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_262_1326 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_17021_ VGND VPWR VGND VPWR _02780_ _02779_ _03145_ keymem.prev_key1_reg\[60\] sky130_fd_sc_hd__a21oi_2
X_14233_ VPWR VGND VGND VPWR _09178_ _09704_ _09091_ sky130_fd_sc_hd__nor2_2
XFILLER_0_227_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_683 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_717 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_22_845 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14164_ VPWR VGND VGND VPWR _09635_ _09633_ _09634_ sky130_fd_sc_hd__nand2_2
XFILLER_0_150_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_150_187 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13115_ VGND VPWR enc_block.round_key\[94\] _08623_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14095_ VGND VPWR VGND VPWR _09353_ _09565_ _09410_ _09441_ _09566_ sky130_fd_sc_hd__o22a_2
X_18972_ VPWR VGND VGND VPWR _04778_ _04806_ _04223_ sky130_fd_sc_hd__nor2_2
XFILLER_0_24_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17923_ VGND VPWR VPWR VGND _03874_ _03879_ keymem.prev_key0_reg\[98\] _03880_ sky130_fd_sc_hd__mux2_2
X_13046_ VPWR VGND VPWR VGND _08560_ keymem.key_mem\[5\]\[88\] _07811_ keymem.key_mem\[8\]\[88\]
+ _07929_ _08561_ sky130_fd_sc_hd__a221o_2
XFILLER_0_237_258 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_219_962 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_158_1507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_206_612 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17854_ VGND VPWR _00217_ _03832_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_238_1553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16805_ VGND VPWR _02866_ key[40] _02949_ _10189_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_234_976 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17785_ VGND VPWR VPWR VGND _03777_ _03096_ keymem.prev_key0_reg\[55\] _03785_ sky130_fd_sc_hd__mux2_2
X_14997_ VPWR VGND VPWR VGND _10424_ _10435_ _10444_ _10419_ _10461_ sky130_fd_sc_hd__or4_2
X_19524_ VGND VPWR VGND VPWR _05162_ keymem.key_mem_we _03119_ _05135_ _00557_ sky130_fd_sc_hd__a31o_2
XFILLER_0_205_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_156_1275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16736_ VPWR VGND VPWR VGND _02886_ keymem.prev_key1_reg\[34\] sky130_fd_sc_hd__inv_2
X_13948_ VGND VPWR VPWR VGND _09328_ _09339_ _09306_ _09420_ sky130_fd_sc_hd__or3_2
XFILLER_0_199_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_92_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19455_ VGND VPWR VGND VPWR _05125_ keymem.key_mem_we _02721_ _05121_ _00525_ sky130_fd_sc_hd__a31o_2
XFILLER_0_5_1001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16667_ VPWR VGND VPWR VGND _02821_ keymem.prev_key0_reg\[126\] sky130_fd_sc_hd__inv_2
X_13879_ VPWR VGND VPWR VGND _09261_ _09317_ _09314_ _09254_ _09351_ sky130_fd_sc_hd__or4_2
XFILLER_0_29_411 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18406_ VPWR VGND VGND VPWR _04297_ _04054_ _04295_ sky130_fd_sc_hd__nand2_2
XFILLER_0_234_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_372 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15618_ VGND VPWR VGND VPWR _11076_ _11075_ _11074_ _10879_ _11073_ sky130_fd_sc_hd__and4_2
XFILLER_0_5_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19386_ VPWR VGND keymem.key_mem_we _05085_ _03654_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16598_ VGND VPWR VGND VPWR _02747_ _02746_ keymem.prev_key1_reg\[123\] _02755_ sky130_fd_sc_hd__a21o_2
XFILLER_0_70_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_45_926 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18337_ VPWR VGND VGND VPWR _04235_ _03961_ _04234_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15549_ VGND VPWR VGND VPWR _10459_ _10482_ _10619_ _10797_ _11008_ sky130_fd_sc_hd__o22a_2
XFILLER_0_44_436 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_112_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18268_ VPWR VGND _04172_ enc_block.block_w2_reg\[10\] enc_block.block_w2_reg\[9\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_245_1513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_114_324 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17219_ VGND VPWR _00091_ _03323_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18199_ VGND VPWR _04109_ enc_block.block_w3_reg\[4\] _04024_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_992 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_163_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20230_ VGND VPWR VPWR VGND _05535_ _09992_ keymem.key_mem\[9\]\[3\] _05539_ sky130_fd_sc_hd__mux2_2
XFILLER_0_124_1219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_177_2_Left_648 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_163_1279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20161_ VGND VPWR _00856_ _05500_ VPWR VGND sky130_fd_sc_hd__buf_1
X_20092_ VGND VPWR _00823_ _05464_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_196_1033 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23920_ VGND VPWR VPWR VGND clk _00413_ reset_n keymem.key_mem\[13\]\[41\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23851_ VGND VPWR VPWR VGND clk _00344_ reset_n enc_block.block_w2_reg\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_240_946 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22802_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[103\] _06858_ _06857_ _05039_ _02139_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_196_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_174_1375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23782_ VGND VPWR VPWR VGND clk _00275_ reset_n enc_block.block_w0_reg\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_71_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20994_ VGND VPWR _01245_ _05944_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_135_1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25521_ VGND VPWR VPWR VGND clk _02014_ reset_n keymem.key_mem\[1\]\[106\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_36_1456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_219 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_22733_ VGND VPWR _02097_ _06831_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_71_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_25452_ VGND VPWR VPWR VGND clk _01945_ reset_n keymem.key_mem\[1\]\[37\] sky130_fd_sc_hd__dfrtp_2
X_22664_ VGND VPWR _02056_ _06803_ VPWR VGND sky130_fd_sc_hd__buf_1
X_21615_ VGND VPWR _01536_ _06274_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24403_ VGND VPWR VPWR VGND clk _00896_ reset_n keymem.key_mem\[9\]\[12\] sky130_fd_sc_hd__dfrtp_2
X_25383_ VGND VPWR VPWR VGND clk _01876_ reset_n keymem.key_mem\[2\]\[96\] sky130_fd_sc_hd__dfrtp_2
X_22595_ VPWR VGND VPWR VGND keymem.key_mem\[1\]\[107\] _06775_ _06774_ _05048_ _02015_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_168_1157 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_164_279 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_24334_ VGND VPWR VPWR VGND clk _00827_ reset_n keymem.key_mem\[10\]\[71\] sky130_fd_sc_hd__dfrtp_2
X_21546_ VGND VPWR VPWR VGND _06231_ _03550_ keymem.key_mem\[5\]\[109\] _06237_ sky130_fd_sc_hd__mux2_2
XFILLER_0_185_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24265_ VGND VPWR VPWR VGND clk _00758_ reset_n keymem.key_mem\[10\]\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_132_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_21477_ VGND VPWR VPWR VGND _06196_ _03295_ keymem.key_mem\[5\]\[76\] _06201_ sky130_fd_sc_hd__mux2_2
X_23216_ VGND VPWR VGND VPWR _07105_ _04266_ _07095_ _07106_ enc_block.block_w3_reg\[1\]
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_120_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_82_1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20428_ VGND VPWR _00981_ _05642_ VPWR VGND sky130_fd_sc_hd__buf_1
X_24196_ VGND VPWR VPWR VGND clk _00689_ reset_n keymem.key_mem\[11\]\[61\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_142_1319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_247_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23147_ VGND VPWR VGND VPWR _03546_ _10085_ _03549_ _07057_ sky130_fd_sc_hd__a21o_2
XFILLER_0_43_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_20359_ VGND VPWR _00948_ _05606_ VPWR VGND sky130_fd_sc_hd__buf_1
X_23078_ VGND VPWR VGND VPWR _06976_ _11555_ _02259_ _07014_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_262_526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_22029_ VGND VPWR VPWR VGND _06494_ _04995_ keymem.key_mem\[3\]\[77\] _06496_ sky130_fd_sc_hd__mux2_2
X_14920_ VPWR VGND _10384_ keymem.prev_key0_reg\[72\] keymem.prev_key0_reg\[40\] VPWR
+ VGND sky130_fd_sc_hd__xor2_2
X_14851_ VPWR VGND _10292_ _10316_ _10315_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_192_1442 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_216_998 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13802_ VPWR VGND VPWR VGND _09274_ enc_block.block_w0_reg\[31\] _09273_ sky130_fd_sc_hd__or2_2
XFILLER_0_187_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_153_1415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_192_1475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17570_ VPWR VGND VPWR VGND _03632_ _03077_ _02733_ _02734_ _03631_ _02496_ sky130_fd_sc_hd__o311a_2
X_14782_ VGND VPWR VPWR VGND _10043_ _10248_ _10247_ sky130_fd_sc_hd__and2b_2
X_11994_ VGND VPWR _07597_ _07596_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_93_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_97_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16521_ VGND VPWR VGND VPWR _02679_ _02678_ _02680_ _02681_ sky130_fd_sc_hd__a21o_2
X_13733_ VGND VPWR VGND VPWR _09129_ _09204_ _09205_ _09141_ sky130_fd_sc_hd__a21oi_2
X_25719_ keymem.prev_key1_reg\[35\] clk _02212_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_50_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19240_ VGND VPWR VPWR VGND _04951_ _04989_ keymem.key_mem\[13\]\[74\] _04990_ sky130_fd_sc_hd__mux2_2
X_16452_ VGND VPWR VPWR VGND _02525_ _02575_ _02519_ _02613_ sky130_fd_sc_hd__or3_2
X_13664_ VGND VPWR _09136_ _09135_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_6_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_112_1145 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_213_40 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15403_ VGND VPWR VGND VPWR _10611_ _10441_ _10455_ _10539_ _10864_ sky130_fd_sc_hd__a31o_2
XFILLER_0_2_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19171_ VGND VPWR _00418_ _04948_ VPWR VGND sky130_fd_sc_hd__buf_1
X_12615_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[45\] _07536_ _08172_ _08168_ _08173_
+ sky130_fd_sc_hd__o22a_2
X_16383_ VGND VPWR VGND VPWR _09717_ _02544_ _02542_ _02543_ _02546_ sky130_fd_sc_hd__a31o_2
X_13595_ VGND VPWR _09067_ _09066_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_213_84 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_155_268 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18122_ VPWR VGND _04039_ _04038_ enc_block.round_key\[101\] VPWR VGND sky130_fd_sc_hd__xor2_2
X_15334_ VGND VPWR VGND VPWR _10513_ _10501_ _10627_ _10530_ _10796_ sky130_fd_sc_hd__o22a_2
XFILLER_0_5_319 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_26_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_1_Right_674 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12546_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[39\] _07562_ keymem.key_mem\[2\]\[39\]
+ _07816_ _08110_ sky130_fd_sc_hd__a22o_2
X_18053_ VGND VPWR VPWR VGND _03974_ enc_block.block_w0_reg\[0\] _03971_ _03975_ sky130_fd_sc_hd__mux2_2
X_15265_ VGND VPWR VGND VPWR _10713_ _10727_ _10728_ _10696_ _10720_ sky130_fd_sc_hd__nor4_2
X_12477_ VPWR VGND VPWR VGND keymem.key_mem\[13\]\[33\] _07812_ keymem.key_mem\[4\]\[33\]
+ _07913_ _08047_ sky130_fd_sc_hd__a22o_2
XFILLER_0_164_1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_491 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_17004_ VGND VPWR _03130_ _03129_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_1_514 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14216_ VGND VPWR _09687_ _09684_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_123_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_160_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15196_ VGND VPWR VGND VPWR _10660_ _10656_ _10385_ _10657_ _10659_ sky130_fd_sc_hd__a211o_2
XFILLER_0_50_973 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_21_152 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_158_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14147_ VPWR VGND VGND VPWR _09410_ _09618_ _09437_ sky130_fd_sc_hd__nor2_2
XFILLER_0_21_174 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_61_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18955_ VPWR VGND _04790_ enc_block.block_w2_reg\[29\] enc_block.block_w3_reg\[20\]
+ VPWR VGND sky130_fd_sc_hd__xor2_2
X_14078_ VPWR VGND VPWR VGND _09549_ _09548_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13029_ VPWR VGND VPWR VGND keymem.key_mem\[7\]\[86\] _08391_ keymem.key_mem\[1\]\[86\]
+ _07670_ _08546_ sky130_fd_sc_hd__a22o_2
X_17906_ VGND VPWR VGND VPWR _03737_ keymem.prev_key1_reg\[93\] _03738_ _03868_ sky130_fd_sc_hd__a21o_2
X_18886_ VPWR VGND VGND VPWR _04728_ enc_block.block_w1_reg\[5\] enc_block.block_w1_reg\[6\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_101_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_17837_ VGND VPWR VPWR VGND _03812_ key[199] keymem.prev_key1_reg\[71\] _03821_ sky130_fd_sc_hd__mux2_2
XFILLER_0_233_250 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_83_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_107_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_171_1515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17768_ VGND VPWR VPWR VGND _03763_ _03032_ keymem.prev_key0_reg\[48\] _03775_ sky130_fd_sc_hd__mux2_2
XFILLER_0_178_327 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16719_ VGND VPWR VGND VPWR keylen _02871_ _02870_ keymem.prev_key1_reg\[32\] _09529_
+ _09530_ sky130_fd_sc_hd__a311oi_2
X_19507_ VGND VPWR _00549_ _05153_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_171_1559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17699_ VGND VPWR _03730_ _03729_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_14_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19438_ VGND VPWR _05116_ _05094_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_18_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_186_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_19369_ VGND VPWR VPWR VGND _05067_ _05073_ keymem.key_mem\[13\]\[119\] _05074_ sky130_fd_sc_hd__mux2_2
X_21400_ VGND VPWR _01435_ _06160_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_84_391 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_242_Left_509 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_22380_ VGND VPWR _01894_ _06681_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_161_238 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_715 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_32_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21331_ VGND VPWR _01402_ _06124_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_5_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_199_66 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_940 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_128_1163 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24050_ VGND VPWR VPWR VGND clk _00543_ reset_n keymem.key_mem\[12\]\[43\] sky130_fd_sc_hd__dfrtp_2
X_21262_ VGND VPWR _01371_ _06086_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_206_1338 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_12_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_12_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23001_ VGND VPWR VGND VPWR _03071_ _03070_ _03074_ _06968_ sky130_fd_sc_hd__a21o_2
XFILLER_0_60_1004 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_20213_ VGND VPWR _00881_ _05527_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_64_1173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_21193_ VGND VPWR _01338_ _06050_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_12_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_40_494 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_556 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_20144_ VGND VPWR _00848_ _05491_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_99_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_217_729 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_251_Left_518 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_24952_ VGND VPWR VPWR VGND clk _01445_ reset_n keymem.key_mem\[5\]\[49\] sky130_fd_sc_hd__dfrtp_2
X_20075_ VGND VPWR _00815_ _05455_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_209_291 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_23903_ VGND VPWR VPWR VGND clk _00396_ reset_n keymem.key_mem\[13\]\[24\] sky130_fd_sc_hd__dfrtp_2
X_24883_ VGND VPWR VPWR VGND clk _01376_ reset_n keymem.key_mem\[6\]\[108\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_217_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1325 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_23834_ VGND VPWR VPWR VGND clk _00327_ reset_n enc_block.block_w1_reg\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_79_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_212_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_135_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1194 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_212_467 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_169_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20977_ VGND VPWR VPWR VGND _05934_ _05027_ keymem.key_mem\[7\]\[97\] _05936_ sky130_fd_sc_hd__mux2_2
X_23765_ keymem.prev_key0_reg\[121\] clk _00262_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_36_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_25504_ VGND VPWR VPWR VGND clk _01997_ reset_n keymem.key_mem\[1\]\[89\] sky130_fd_sc_hd__dfrtp_2
X_22716_ VPWR VGND VPWR VGND keymem.key_mem\[0\]\[52\] _06820_ _06819_ _04958_ _02088_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_3_1505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_23696_ keymem.prev_key0_reg\[52\] clk _00193_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_250_1093 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_36_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_71_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_260_Left_527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_25435_ VGND VPWR VPWR VGND clk _01928_ reset_n keymem.key_mem\[1\]\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_1549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_22647_ VGND VPWR _02048_ _06794_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_75_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12400_ VPWR VGND VPWR VGND _07976_ keymem.key_mem\[9\]\[26\] _07612_ keymem.key_mem\[8\]\[26\]
+ _07903_ _07977_ sky130_fd_sc_hd__a221o_2
XFILLER_0_24_907 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13380_ VPWR VGND VPWR VGND keymem.key_mem\[10\]\[121\] _07562_ keymem.key_mem\[1\]\[121\]
+ _07558_ _08862_ sky130_fd_sc_hd__a22o_2
X_25366_ VGND VPWR VPWR VGND clk _01859_ reset_n keymem.key_mem\[2\]\[79\] sky130_fd_sc_hd__dfrtp_2
X_22578_ VGND VPWR _02001_ _06772_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_228_1541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24317_ VGND VPWR VPWR VGND clk _00810_ reset_n keymem.key_mem\[10\]\[54\] sky130_fd_sc_hd__dfrtp_2
X_12331_ VGND VPWR _07914_ _07913_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_1_1284 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_63_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21529_ VGND VPWR VPWR VGND _06220_ _03499_ keymem.key_mem\[5\]\[101\] _06228_ sky130_fd_sc_hd__mux2_2
X_25297_ VGND VPWR VPWR VGND clk _01790_ reset_n keymem.key_mem\[2\]\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_105_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15050_ VGND VPWR _10514_ _10451_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_32_951 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12262_ VPWR VGND VPWR VGND keymem.key_mem\[11\]\[15\] _07631_ keymem.key_mem\[2\]\[15\]
+ _07697_ _07850_ sky130_fd_sc_hd__a22o_2
XFILLER_0_146_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24248_ VGND VPWR VPWR VGND clk _00741_ reset_n keymem.key_mem\[11\]\[113\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_267_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14001_ VPWR VGND VGND VPWR _09341_ _09473_ _09303_ sky130_fd_sc_hd__nor2_2
XFILLER_0_107_1247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_259_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_472 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_483 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_24179_ VGND VPWR VPWR VGND clk _00672_ reset_n keymem.key_mem\[11\]\[44\] sky130_fd_sc_hd__dfrtp_2
X_12193_ VGND VPWR _07786_ _07785_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_82_1295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_208_718 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_247_364 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_101_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_128_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18740_ _04594_ _04596_ _04065_ _04595_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_37_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15952_ VGND VPWR VGND VPWR _11408_ _11273_ _11228_ _11272_ _11226_ sky130_fd_sc_hd__and4_2
XFILLER_0_235_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_740 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_262_356 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14903_ VPWR VGND VGND VPWR _10368_ _10367_ _10365_ _10328_ _10327_ key[7] sky130_fd_sc_hd__o2111a_2
X_18671_ VPWR VGND VGND VPWR _04512_ _04535_ _04240_ sky130_fd_sc_hd__nor2_2
XFILLER_0_204_902 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15883_ VGND VPWR VGND VPWR _11339_ _11273_ _11289_ _11272_ _11226_ sky130_fd_sc_hd__and4_2
X_17622_ VGND VPWR _00141_ _03676_ VPWR VGND sky130_fd_sc_hd__buf_1
X_14834_ VGND VPWR VGND VPWR _10299_ _10297_ _09401_ _09333_ _10298_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_53_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_187_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_303 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_114_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17553_ VGND VPWR VGND VPWR _02679_ _02678_ _03617_ _10967_ sky130_fd_sc_hd__a21oi_2
X_14765_ VPWR VGND VPWR VGND _09550_ _09553_ _09360_ _09464_ _10231_ sky130_fd_sc_hd__a22o_2
XFILLER_0_93_1391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11977_ VGND VPWR _07580_ _07579_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_212_990 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_16504_ VGND VPWR VGND VPWR keymem.rcon_reg\[0\] _11301_ _02664_ _11438_ sky130_fd_sc_hd__a21bo_2
X_13716_ VGND VPWR VGND VPWR _09188_ _09015_ _08991_ _09014_ _09043_ sky130_fd_sc_hd__and4_2
XFILLER_0_15_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_17484_ VGND VPWR VGND VPWR _03557_ _03302_ _08937_ key[111] sky130_fd_sc_hd__o21a_2
X_14696_ VGND VPWR VGND VPWR _09136_ _09113_ _09153_ _09125_ _10163_ sky130_fd_sc_hd__o22a_2
XFILLER_0_54_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19223_ VPWR VGND keymem.key_mem\[13\]\[67\] _04980_ _04979_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_6_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16435_ VGND VPWR keymem.prev_key1_reg\[118\] _11072_ _02597_ _11089_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_13647_ VPWR VGND VGND VPWR _09119_ _09104_ _09118_ sky130_fd_sc_hd__nand2_2
XFILLER_0_160_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_606 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_85_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_363 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_128_279 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_19154_ VPWR VGND keymem.key_mem_we _04937_ _02964_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_6_639 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_16366_ VPWR VGND VGND VPWR _02528_ _02527_ _11323_ _11389_ _11434_ _02529_ sky130_fd_sc_hd__a311o_2
XFILLER_0_27_778 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13578_ VGND VPWR _09050_ _09049_ VPWR VGND sky130_fd_sc_hd__buf_1
X_18105_ VPWR VGND _04023_ _04022_ _04021_ VPWR VGND sky130_fd_sc_hd__xor2_2
X_15317_ VGND VPWR VGND VPWR _10462_ _10497_ _10557_ _10503_ _10779_ sky130_fd_sc_hd__o22a_2
XPHY_EDGE_ROW_74_1_Right_675 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12529_ VGND VPWR VGND VPWR keymem.key_mem\[0\]\[37\] _07893_ _08094_ _08089_ _08095_
+ sky130_fd_sc_hd__o22a_2
X_19085_ VPWR VGND keymem.key_mem\[13\]\[12\] _04897_ _04887_ VPWR VGND sky130_fd_sc_hd__and2_2
X_16297_ VGND VPWR VGND VPWR _02459_ keymem.prev_key0_reg\[116\] _02461_ _02412_ sky130_fd_sc_hd__nand3_2
XFILLER_0_240_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18036_ VGND VPWR _03958_ _03957_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_125_1303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15248_ VGND VPWR VGND VPWR _10584_ _10604_ _10475_ _10458_ _10553_ _10711_ sky130_fd_sc_hd__o32a_2
XFILLER_0_78_23 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_164_1363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_65_1471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_125_1347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_355 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15179_ VGND VPWR VGND VPWR _10638_ _10472_ _10640_ _10641_ _10643_ _10642_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_10_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_254_802 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_238_353 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_254_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_19987_ VGND VPWR _00773_ _05409_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_185_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_18938_ VPWR VGND VGND VPWR _04774_ _04775_ _04478_ sky130_fd_sc_hd__nor2_2
XFILLER_0_185_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
.ends

