../007-success-hybrid-abstract-gds/spm.lef